library IEEE;
use IEEE.std_logic_1164.all;

--  A testbench has no ports.
entity dregister_tb is
end dregister_tb;

architecture dregister_tb_arch of dregister_tb is
   --  Declaration of the component that will be instantiated.
   component dregister
     port (d : in std_logic_vector(15 downto 0); load, clk : in std_logic; cout : out std_logic_vector(15 downto 0));
   end component;
   -- Declaration of the clock
   component Clock
     port (finish : in std_logic;
           cout   : out std_logic);
   end component;
   
   --  Specifies which entity is bound with the component.
   for dregister_0: dregister use entity work.dregister;
   signal d, cout : std_logic_vector(15 downto 0);
   signal load, finish, clk : std_logic;
begin
  --  Component instantiation.
  OSC_CLK: Clock port map (finish, clk);
  dregister_0: dregister port map (d, load, clk, cout);

   --  This process does the real job.
   process
      type pattern_type is record
         --  The inputs of the dregister.
        d    : std_logic_vector(15 downto 0);
        load : std_logic;
        --  The output of the dregister.
        cout : std_logic_vector(15 downto 0);
      end record;
      --  The patterns to apply.
      type pattern_array is array (natural range <>) of pattern_type;
      constant patterns : pattern_array :=
        (("0000000000000000", '0', "0000000000000000"),
         ("0000000000000000", '0', "0000000000000000"),
         ("0000000000000000", '1', "0000000000000000"),
         ("0000000000000000", '1', "0000000000000000"),
         ("0111110101111011", '0', "0000000000000000"),
         ("0111110101111011", '0', "0000000000000000"),
         ("0010101101100111", '0', "0000000000000000"),
         ("0010101101100111", '0', "0000000000000000"),
         ("0111110101111011", '1', "0000000000000000"),
         ("0111110101111011", '1', "0111110101111011"),
         ("0111110101111011", '1', "0111110101111011"),
         ("0111110101111011", '1', "0111110101111011"),
         ("0111110101111011", '0', "0111110101111011"),
         ("0111110101111011", '0', "0111110101111011"),
         ("0011000000111001", '1', "0111110101111011"),
         ("0011000000111001", '1', "0011000000111001"),
         ("0000000000000000", '0', "0011000000111001"),
         ("0000000000000000", '0', "0011000000111001"),
         ("0000000000000000", '1', "0011000000111001"),
         ("0000000000000000", '1', "0000000000000000"),
         ("0000000000000001", '0', "0000000000000000"),
         ("0000000000000001", '0', "0000000000000000"),
         ("0000000000000001", '1', "0000000000000000"),
         ("0000000000000001", '1', "0000000000000001"),
         ("0000000000000010", '0', "0000000000000001"),
         ("0000000000000010", '0', "0000000000000001"),
         ("0000000000000010", '1', "0000000000000001"),
         ("0000000000000010", '1', "0000000000000010"),
         ("0000000000000100", '0', "0000000000000010"),
         ("0000000000000100", '0', "0000000000000010"),
         ("0000000000000100", '1', "0000000000000010"),
         ("0000000000000100", '1', "0000000000000100"),
         ("0000000000001000", '0', "0000000000000100"),
         ("0000000000001000", '0', "0000000000000100"),
         ("0000000000001000", '1', "0000000000000100"),
         ("0000000000001000", '1', "0000000000001000"),
         ("0000000000010000", '0', "0000000000001000"),
         ("0000000000010000", '0', "0000000000001000"),
         ("0000000000010000", '1', "0000000000001000"),
         ("0000000000010000", '1', "0000000000010000"),
         ("0000000000100000", '0', "0000000000010000"),
         ("0000000000100000", '0', "0000000000010000"),
         ("0000000000100000", '1', "0000000000010000"),
         ("0000000000100000", '1', "0000000000100000"),
         ("0000000001000000", '0', "0000000000100000"),
         ("0000000001000000", '0', "0000000000100000"),
         ("0000000001000000", '1', "0000000000100000"),
         ("0000000001000000", '1', "0000000001000000"),
         ("0000000010000000", '0', "0000000001000000"),
         ("0000000010000000", '0', "0000000001000000"),
         ("0000000010000000", '1', "0000000001000000"),
         ("0000000010000000", '1', "0000000010000000"),
         ("0000000100000000", '0', "0000000010000000"),
         ("0000000100000000", '0', "0000000010000000"),
         ("0000000100000000", '1', "0000000010000000"),
         ("0000000100000000", '1', "0000000100000000"),
         ("0000001000000000", '0', "0000000100000000"),
         ("0000001000000000", '0', "0000000100000000"),
         ("0000001000000000", '1', "0000000100000000"),
         ("0000001000000000", '1', "0000001000000000"),
         ("0000010000000000", '0', "0000001000000000"),
         ("0000010000000000", '0', "0000001000000000"),
         ("0000010000000000", '1', "0000001000000000"),
         ("0000010000000000", '1', "0000010000000000"),
         ("0000100000000000", '0', "0000010000000000"),
         ("0000100000000000", '0', "0000010000000000"),
         ("0000100000000000", '1', "0000010000000000"),
         ("0000100000000000", '1', "0000100000000000"),
         ("0001000000000000", '0', "0000100000000000"),
         ("0001000000000000", '0', "0000100000000000"),
         ("0001000000000000", '1', "0000100000000000"),
         ("0001000000000000", '1', "0001000000000000"),
         ("0010000000000000", '0', "0001000000000000"),
         ("0010000000000000", '0', "0001000000000000"),
         ("0010000000000000", '1', "0001000000000000"),
         ("0010000000000000", '1', "0010000000000000"),
         ("0100000000000000", '0', "0010000000000000"),
         ("0100000000000000", '0', "0010000000000000"),
         ("0100000000000000", '1', "0010000000000000"),
         ("0100000000000000", '1', "0100000000000000"),
         ("1000000000000000", '0', "0100000000000000"),
         ("1000000000000000", '0', "0100000000000000"),
         ("1000000000000000", '1', "0100000000000000"),
         ("1000000000000000", '1', "1000000000000000"),
         ("0000000000000010", '0', "1000000000000000"),
         ("0000000000000010", '0', "1000000000000000"),
         ("0000000000000010", '1', "1000000000000000"),
         ("0000000000000010", '1', "0000000000000010"),
         ("0000000000000011", '0', "0000000000000010"),
         ("0000000000000011", '0', "0000000000000010"),
         ("0000000000000011", '1', "0000000000000010"),
         ("0000000000000011", '1', "0000000000000011"),
         ("0000000000000101", '0', "0000000000000011"),
         ("0000000000000101", '0', "0000000000000011"),
         ("0000000000000101", '1', "0000000000000011"),
         ("0000000000000101", '1', "0000000000000101"),
         ("0000000000001001", '0', "0000000000000101"),
         ("0000000000001001", '0', "0000000000000101"),
         ("0000000000001001", '1', "0000000000000101"),
         ("0000000000001001", '1', "0000000000001001"),
         ("0000000000010001", '0', "0000000000001001"),
         ("0000000000010001", '0', "0000000000001001"),
         ("0000000000010001", '1', "0000000000001001"),
         ("0000000000010001", '1', "0000000000010001"),
         ("0000000000100001", '0', "0000000000010001"),
         ("0000000000100001", '0', "0000000000010001"),
         ("0000000000100001", '1', "0000000000010001"),
         ("0000000000100001", '1', "0000000000100001"),
         ("0000000001000001", '0', "0000000000100001"),
         ("0000000001000001", '0', "0000000000100001"),
         ("0000000001000001", '1', "0000000000100001"),
         ("0000000001000001", '1', "0000000001000001"),
         ("0000000010000001", '0', "0000000001000001"),
         ("0000000010000001", '0', "0000000001000001"),
         ("0000000010000001", '1', "0000000001000001"),
         ("0000000010000001", '1', "0000000010000001"),
         ("0000000100000001", '0', "0000000010000001"),
         ("0000000100000001", '0', "0000000010000001"),
         ("0000000100000001", '1', "0000000010000001"),
         ("0000000100000001", '1', "0000000100000001"),
         ("0000001000000001", '0', "0000000100000001"),
         ("0000001000000001", '0', "0000000100000001"),
         ("0000001000000001", '1', "0000000100000001"),
         ("0000001000000001", '1', "0000001000000001"),
         ("0000010000000001", '0', "0000001000000001"),
         ("0000010000000001", '0', "0000001000000001"),
         ("0000010000000001", '1', "0000001000000001"),
         ("0000010000000001", '1', "0000010000000001"),
         ("0000100000000001", '0', "0000010000000001"),
         ("0000100000000001", '0', "0000010000000001"),
         ("0000100000000001", '1', "0000010000000001"),
         ("0000100000000001", '1', "0000100000000001"),
         ("0001000000000001", '0', "0000100000000001"),
         ("0001000000000001", '0', "0000100000000001"),
         ("0001000000000001", '1', "0000100000000001"),
         ("0001000000000001", '1', "0001000000000001"),
         ("0010000000000001", '0', "0001000000000001"),
         ("0010000000000001", '0', "0001000000000001"),
         ("0010000000000001", '1', "0001000000000001"),
         ("0010000000000001", '1', "0010000000000001"),
         ("0100000000000001", '0', "0010000000000001"),
         ("0100000000000001", '0', "0010000000000001"),
         ("0100000000000001", '1', "0010000000000001"),
         ("0100000000000001", '1', "0100000000000001"),
         ("0111111111111111", '0', "0100000000000001"),
         ("0111111111111111", '0', "0100000000000001"),
         ("0111111111111111", '1', "0100000000000001"),
         ("0111111111111111", '1', "0111111111111111"));
         
   begin
      --  Check each pattern.
      for i in patterns'range loop
         --  Set the inputs.
        d <= patterns(i).d;
        load <= patterns(i).load;
        wait for 0.25 ns;
        --  Check the outputs.
        assert cout = patterns(i).cout
          report "bad data; nothing remembered" severity error;
        wait for 0.75 ns;
     end loop;
     -- End the clock
     finish <= '1';
     assert false report "end of test" severity note;
     --  Wait forever; this will finish the simulation.
     wait;
  end process;
end dregister_tb_arch;
