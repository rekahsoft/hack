library IEEE;
use IEEE.std_logic_1164.all;

--  A testbench has no ports.
entity ram16k_tb is
end ram16k_tb;

architecture ram16k_tb_arch of ram16k_tb is
   --  Declaration of the component that will be instantiated.
   component ram16k
     port (d       : in std_logic_vector(15 downto 0);
           load    : in std_logic;
           address : in std_logic_vector(14 downto 0);
           clk     : in std_logic;
           cout    : out std_logic_vector(15 downto 0));
   end component;
   -- Declaration of the clock
   component Clock
     port (finish : in std_logic;
           cout   : out std_logic);
   end component;
   
   --  Specifies which entity is bound with the component.
   for ram16k_0: ram16k use entity work.ram16k;
   signal d, cout : std_logic_vector(15 downto 0);
   signal address : std_logic_vector(14 downto 0);
   signal load, finish, clk : std_logic;
begin
  --  Component instantiation.
  OSC_CLK: Clock port map (finish, clk);
  ram16k_0: ram16k port map (d, load, address, clk, cout);

   --  This process does the real job.
   process
      type pattern_type is record
         --  The inputs of the ram16k.
        d       : std_logic_vector(15 downto 0);
        load    : std_logic;
        address : std_logic_vector(14 downto 0);
        --  The output of the ram16k.
        cout    : std_logic_vector(15 downto 0);
      end record;
      --  The patterns to apply.
      type pattern_array is array (natural range <>) of pattern_type;
      constant patterns : pattern_array :=
        (("0000000000000000", '0', "000000000000000", "0000000000000000"),
         ("0000000000000000", '0', "000000000000000", "0000000000000000"),
         ("0000000000000000", '1', "000000000000000", "0000000000000000"),
         ("0000000000000000", '1', "000000000000000", "0000000000000000"),
         ("0001000011100001", '0', "000000000000000", "0000000000000000"),
         ("0001000011100001", '0', "000000000000000", "0000000000000000"),
         ("0001000011100001", '1', "001000011100001", "0000000000000000"),
         ("0001000011100001", '1', "001000011100001", "0001000011100001"),
         ("0001000011100001", '0', "000000000000000", "0000000000000000"),
         ("0001000011100001", '0', "000000000000000", "0000000000000000"),
         ("0011000000111001", '0', "011000000111001", "0000000000000000"),
         ("0011000000111001", '0', "011000000111001", "0000000000000000"),
         ("0011000000111001", '1', "011000000111001", "0000000000000000"),
         ("0011000000111001", '1', "011000000111001", "0011000000111001"),
         ("0011000000111001", '0', "011000000111001", "0011000000111001"),
         ("0011000000111001", '0', "011000000111001", "0011000000111001"),
         ("0011000000111001", '0', "001000011100001", "0001000011100001"),
         ("0011111111111111", '0', "001000011100001", "0001000011100001"),
         ("0011111111111111", '0', "001000011100001", "0001000011100001"),
         ("0011111111111111", '1', "011111111111111", "0000000000000000"),
         ("0011111111111111", '1', "011111111111111", "0011111111111111"),
         ("0011111111111111", '0', "011111111111111", "0011111111111111"),
         ("0011111111111111", '0', "011111111111111", "0011111111111111"),
         ("0011111111111111", '0', "011000000111001", "0011000000111001"),
         ("0011111111111111", '0', "011111111111111", "0011111111111111"),
         ("0011111111111111", '0', "010101010101000", "0000000000000000"),
         ("0011111111111111", '0', "010101010101000", "0000000000000000"),
         ("0011111111111111", '0', "010101010101001", "0000000000000000"),
         ("0011111111111111", '0', "010101010101010", "0000000000000000"),
         ("0011111111111111", '0', "010101010101011", "0000000000000000"),
         ("0011111111111111", '0', "010101010101100", "0000000000000000"),
         ("0011111111111111", '0', "010101010101101", "0000000000000000"),
         ("0011111111111111", '0', "010101010101110", "0000000000000000"),
         ("0011111111111111", '0', "010101010101111", "0000000000000000"),
         ("0101010101010101", '1', "010101010101000", "0000000000000000"),
         ("0101010101010101", '1', "010101010101000", "0101010101010101"),
         ("0101010101010101", '1', "010101010101001", "0000000000000000"),
         ("0101010101010101", '1', "010101010101001", "0101010101010101"),
         ("0101010101010101", '1', "010101010101010", "0000000000000000"),
         ("0101010101010101", '1', "010101010101010", "0101010101010101"),
         ("0101010101010101", '1', "010101010101011", "0000000000000000"),
         ("0101010101010101", '1', "010101010101011", "0101010101010101"),
         ("0101010101010101", '1', "010101010101100", "0000000000000000"),
         ("0101010101010101", '1', "010101010101100", "0101010101010101"),
         ("0101010101010101", '1', "010101010101101", "0000000000000000"),
         ("0101010101010101", '1', "010101010101101", "0101010101010101"),
         ("0101010101010101", '1', "010101010101110", "0000000000000000"),
         ("0101010101010101", '1', "010101010101110", "0101010101010101"),
         ("0101010101010101", '1', "010101010101111", "0000000000000000"),
         ("0101010101010101", '1', "010101010101111", "0101010101010101"),
         ("0101010101010101", '0', "010101010101000", "0101010101010101"),
         ("0101010101010101", '0', "010101010101000", "0101010101010101"),
         ("0101010101010101", '0', "010101010101001", "0101010101010101"),
         ("0101010101010101", '0', "010101010101010", "0101010101010101"),
         ("0101010101010101", '0', "010101010101011", "0101010101010101"),
         ("0101010101010101", '0', "010101010101100", "0101010101010101"),
         ("0101010101010101", '0', "010101010101101", "0101010101010101"),
         ("0101010101010101", '0', "010101010101110", "0101010101010101"),
         ("0101010101010101", '0', "010101010101111", "0101010101010101"),
         ("0101010101010110", '1', "010101010101000", "0101010101010101"),
         ("0101010101010110", '1', "010101010101000", "0101010101010110"),
         ("0101010101010110", '0', "010101010101000", "0101010101010110"),
         ("0101010101010110", '0', "010101010101000", "0101010101010110"),
         ("0101010101010110", '0', "010101010101001", "0101010101010101"),
         ("0101010101010110", '0', "010101010101010", "0101010101010101"),
         ("0101010101010110", '0', "010101010101011", "0101010101010101"),
         ("0101010101010110", '0', "010101010101100", "0101010101010101"),
         ("0101010101010110", '0', "010101010101101", "0101010101010101"),
         ("0101010101010110", '0', "010101010101110", "0101010101010101"),
         ("0101010101010110", '0', "010101010101111", "0101010101010101"),
         ("0101010101010101", '1', "010101010101000", "0101010101010110"),
         ("0101010101010101", '1', "010101010101000", "0101010101010101"),
         ("0101010101010110", '1', "010101010101001", "0101010101010101"),
         ("0101010101010110", '1', "010101010101001", "0101010101010110"),
         ("0101010101010110", '0', "010101010101000", "0101010101010101"),
         ("0101010101010110", '0', "010101010101000", "0101010101010101"),
         ("0101010101010110", '0', "010101010101001", "0101010101010110"),
         ("0101010101010110", '0', "010101010101010", "0101010101010101"),
         ("0101010101010110", '0', "010101010101011", "0101010101010101"),
         ("0101010101010110", '0', "010101010101100", "0101010101010101"),
         ("0101010101010110", '0', "010101010101101", "0101010101010101"),
         ("0101010101010110", '0', "010101010101110", "0101010101010101"),
         ("0101010101010110", '0', "010101010101111", "0101010101010101"),
         ("0101010101010101", '1', "010101010101001", "0101010101010110"),
         ("0101010101010101", '1', "010101010101001", "0101010101010101"),
         ("0101010101010110", '1', "010101010101010", "0101010101010101"),
         ("0101010101010110", '1', "010101010101010", "0101010101010110"),
         ("0101010101010110", '0', "010101010101000", "0101010101010101"),
         ("0101010101010110", '0', "010101010101000", "0101010101010101"),
         ("0101010101010110", '0', "010101010101001", "0101010101010101"),
         ("0101010101010110", '0', "010101010101010", "0101010101010110"),
         ("0101010101010110", '0', "010101010101011", "0101010101010101"),
         ("0101010101010110", '0', "010101010101100", "0101010101010101"),
         ("0101010101010110", '0', "010101010101101", "0101010101010101"),
         ("0101010101010110", '0', "010101010101110", "0101010101010101"),
         ("0101010101010110", '0', "010101010101111", "0101010101010101"),
         ("0101010101010101", '1', "010101010101010", "0101010101010110"),
         ("0101010101010101", '1', "010101010101010", "0101010101010101"),
         ("0101010101010110", '1', "010101010101011", "0101010101010101"),
         ("0101010101010110", '1', "010101010101011", "0101010101010110"),
         ("0101010101010110", '0', "010101010101000", "0101010101010101"),
         ("0101010101010110", '0', "010101010101000", "0101010101010101"),
         ("0101010101010110", '0', "010101010101001", "0101010101010101"),
         ("0101010101010110", '0', "010101010101010", "0101010101010101"),
         ("0101010101010110", '0', "010101010101011", "0101010101010110"),
         ("0101010101010110", '0', "010101010101100", "0101010101010101"),
         ("0101010101010110", '0', "010101010101101", "0101010101010101"),
         ("0101010101010110", '0', "010101010101110", "0101010101010101"),
         ("0101010101010110", '0', "010101010101111", "0101010101010101"),
         ("0101010101010101", '1', "010101010101011", "0101010101010110"),
         ("0101010101010101", '1', "010101010101011", "0101010101010101"),
         ("0101010101010110", '1', "010101010101100", "0101010101010101"),
         ("0101010101010110", '1', "010101010101100", "0101010101010110"),
         ("0101010101010110", '0', "010101010101000", "0101010101010101"),
         ("0101010101010110", '0', "010101010101000", "0101010101010101"),
         ("0101010101010110", '0', "010101010101001", "0101010101010101"),
         ("0101010101010110", '0', "010101010101010", "0101010101010101"),
         ("0101010101010110", '0', "010101010101011", "0101010101010101"),
         ("0101010101010110", '0', "010101010101100", "0101010101010110"),
         ("0101010101010110", '0', "010101010101101", "0101010101010101"),
         ("0101010101010110", '0', "010101010101110", "0101010101010101"),
         ("0101010101010110", '0', "010101010101111", "0101010101010101"),
         ("0101010101010101", '1', "010101010101100", "0101010101010110"),
         ("0101010101010101", '1', "010101010101100", "0101010101010101"),
         ("0101010101010110", '1', "010101010101101", "0101010101010101"),
         ("0101010101010110", '1', "010101010101101", "0101010101010110"),
         ("0101010101010110", '0', "010101010101000", "0101010101010101"),
         ("0101010101010110", '0', "010101010101000", "0101010101010101"),
         ("0101010101010110", '0', "010101010101001", "0101010101010101"),
         ("0101010101010110", '0', "010101010101010", "0101010101010101"),
         ("0101010101010110", '0', "010101010101011", "0101010101010101"),
         ("0101010101010110", '0', "010101010101100", "0101010101010101"),
         ("0101010101010110", '0', "010101010101101", "0101010101010110"),
         ("0101010101010110", '0', "010101010101110", "0101010101010101"),
         ("0101010101010110", '0', "010101010101111", "0101010101010101"),
         ("0101010101010101", '1', "010101010101101", "0101010101010110"),
         ("0101010101010101", '1', "010101010101101", "0101010101010101"),
         ("0101010101010110", '1', "010101010101110", "0101010101010101"),
         ("0101010101010110", '1', "010101010101110", "0101010101010110"),
         ("0101010101010110", '0', "010101010101000", "0101010101010101"),
         ("0101010101010110", '0', "010101010101000", "0101010101010101"),
         ("0101010101010110", '0', "010101010101001", "0101010101010101"),
         ("0101010101010110", '0', "010101010101010", "0101010101010101"),
         ("0101010101010110", '0', "010101010101011", "0101010101010101"),
         ("0101010101010110", '0', "010101010101100", "0101010101010101"),
         ("0101010101010110", '0', "010101010101101", "0101010101010101"),
         ("0101010101010110", '0', "010101010101110", "0101010101010110"),
         ("0101010101010110", '0', "010101010101111", "0101010101010101"),
         ("0101010101010101", '1', "010101010101110", "0101010101010110"),
         ("0101010101010101", '1', "010101010101110", "0101010101010101"),
         ("0101010101010110", '1', "010101010101111", "0101010101010101"),
         ("0101010101010110", '1', "010101010101111", "0101010101010110"),
         ("0101010101010110", '0', "010101010101000", "0101010101010101"),
         ("0101010101010110", '0', "010101010101000", "0101010101010101"),
         ("0101010101010110", '0', "010101010101001", "0101010101010101"),
         ("0101010101010110", '0', "010101010101010", "0101010101010101"),
         ("0101010101010110", '0', "010101010101011", "0101010101010101"),
         ("0101010101010110", '0', "010101010101100", "0101010101010101"),
         ("0101010101010110", '0', "010101010101101", "0101010101010101"),
         ("0101010101010110", '0', "010101010101110", "0101010101010101"),
         ("0101010101010110", '0', "010101010101111", "0101010101010110"),
         ("0101010101010101", '1', "010101010101111", "0101010101010110"),
         ("0101010101010101", '1', "010101010101111", "0101010101010101"),
         ("0101010101010101", '0', "010101010101000", "0101010101010101"),
         ("0101010101010101", '0', "010101010101000", "0101010101010101"),
         ("0101010101010101", '0', "010101010101001", "0101010101010101"),
         ("0101010101010101", '0', "010101010101010", "0101010101010101"),
         ("0101010101010101", '0', "010101010101011", "0101010101010101"),
         ("0101010101010101", '0', "010101010101100", "0101010101010101"),
         ("0101010101010101", '0', "010101010101101", "0101010101010101"),
         ("0101010101010101", '0', "010101010101110", "0101010101010101"),
         ("0101010101010101", '0', "010101010101111", "0101010101010101"),
         ("0101010101010101", '0', "000010101010101", "0000000000000000"),
         ("0101010101010101", '0', "000010101010101", "0000000000000000"),
         ("0101010101010101", '0', "000110101010101", "0000000000000000"),
         ("0101010101010101", '0', "001010101010101", "0000000000000000"),
         ("0101010101010101", '0', "001110101010101", "0000000000000000"),
         ("0101010101010101", '0', "010010101010101", "0000000000000000"),
         ("0101010101010101", '0', "010110101010101", "0000000000000000"),
         ("0101010101010101", '0', "011010101010101", "0000000000000000"),
         ("0101010101010101", '0', "011110101010101", "0000000000000000"),
         ("0101010101010101", '1', "000010101010101", "0000000000000000"),
         ("0101010101010101", '1', "000010101010101", "0101010101010101"),
         ("0101010101010101", '1', "000110101010101", "0000000000000000"),
         ("0101010101010101", '1', "000110101010101", "0101010101010101"),
         ("0101010101010101", '1', "001010101010101", "0000000000000000"),
         ("0101010101010101", '1', "001010101010101", "0101010101010101"),
         ("0101010101010101", '1', "001110101010101", "0000000000000000"),
         ("0101010101010101", '1', "001110101010101", "0101010101010101"),
         ("0101010101010101", '1', "010010101010101", "0000000000000000"),
         ("0101010101010101", '1', "010010101010101", "0101010101010101"),
         ("0101010101010101", '1', "010110101010101", "0000000000000000"),
         ("0101010101010101", '1', "010110101010101", "0101010101010101"),
         ("0101010101010101", '1', "011010101010101", "0000000000000000"),
         ("0101010101010101", '1', "011010101010101", "0101010101010101"),
         ("0101010101010101", '1', "011110101010101", "0000000000000000"),
         ("0101010101010101", '1', "011110101010101", "0101010101010101"),
         ("0101010101010101", '0', "000010101010101", "0101010101010101"),
         ("0101010101010101", '0', "000010101010101", "0101010101010101"),
         ("0101010101010101", '0', "000110101010101", "0101010101010101"),
         ("0101010101010101", '0', "001010101010101", "0101010101010101"),
         ("0101010101010101", '0', "001110101010101", "0101010101010101"),
         ("0101010101010101", '0', "010010101010101", "0101010101010101"),
         ("0101010101010101", '0', "010110101010101", "0101010101010101"),
         ("0101010101010101", '0', "011010101010101", "0101010101010101"),
         ("0101010101010101", '0', "011110101010101", "0101010101010101"),
         ("0101010101010110", '1', "000010101010101", "0101010101010101"),
         ("0101010101010110", '1', "000010101010101", "0101010101010110"),
         ("0101010101010110", '0', "000010101010101", "0101010101010110"),
         ("0101010101010110", '0', "000010101010101", "0101010101010110"),
         ("0101010101010110", '0', "000110101010101", "0101010101010101"),
         ("0101010101010110", '0', "001010101010101", "0101010101010101"),
         ("0101010101010110", '0', "001110101010101", "0101010101010101"),
         ("0101010101010110", '0', "010010101010101", "0101010101010101"),
         ("0101010101010110", '0', "010110101010101", "0101010101010101"),
         ("0101010101010110", '0', "011010101010101", "0101010101010101"),
         ("0101010101010110", '0', "011110101010101", "0101010101010101"),
         ("0101010101010101", '1', "000010101010101", "0101010101010110"),
         ("0101010101010101", '1', "000010101010101", "0101010101010101"),
         ("0101010101010110", '1', "000110101010101", "0101010101010101"),
         ("0101010101010110", '1', "000110101010101", "0101010101010110"),
         ("0101010101010110", '0', "000010101010101", "0101010101010101"),
         ("0101010101010110", '0', "000010101010101", "0101010101010101"),
         ("0101010101010110", '0', "000110101010101", "0101010101010110"),
         ("0101010101010110", '0', "001010101010101", "0101010101010101"),
         ("0101010101010110", '0', "001110101010101", "0101010101010101"),
         ("0101010101010110", '0', "010010101010101", "0101010101010101"),
         ("0101010101010110", '0', "010110101010101", "0101010101010101"),
         ("0101010101010110", '0', "011010101010101", "0101010101010101"),
         ("0101010101010110", '0', "011110101010101", "0101010101010101"),
         ("0101010101010101", '1', "000110101010101", "0101010101010110"),
         ("0101010101010101", '1', "000110101010101", "0101010101010101"),
         ("0101010101010110", '1', "001010101010101", "0101010101010101"),
         ("0101010101010110", '1', "001010101010101", "0101010101010110"),
         ("0101010101010110", '0', "000010101010101", "0101010101010101"),
         ("0101010101010110", '0', "000010101010101", "0101010101010101"),
         ("0101010101010110", '0', "000110101010101", "0101010101010101"),
         ("0101010101010110", '0', "001010101010101", "0101010101010110"),
         ("0101010101010110", '0', "001110101010101", "0101010101010101"),
         ("0101010101010110", '0', "010010101010101", "0101010101010101"),
         ("0101010101010110", '0', "010110101010101", "0101010101010101"),
         ("0101010101010110", '0', "011010101010101", "0101010101010101"),
         ("0101010101010110", '0', "011110101010101", "0101010101010101"),
         ("0101010101010101", '1', "001010101010101", "0101010101010110"),
         ("0101010101010101", '1', "001010101010101", "0101010101010101"),
         ("0101010101010110", '1', "001110101010101", "0101010101010101"),
         ("0101010101010110", '1', "001110101010101", "0101010101010110"),
         ("0101010101010110", '0', "000010101010101", "0101010101010101"),
         ("0101010101010110", '0', "000010101010101", "0101010101010101"),
         ("0101010101010110", '0', "000110101010101", "0101010101010101"),
         ("0101010101010110", '0', "001010101010101", "0101010101010101"),
         ("0101010101010110", '0', "001110101010101", "0101010101010110"),
         ("0101010101010110", '0', "010010101010101", "0101010101010101"),
         ("0101010101010110", '0', "010110101010101", "0101010101010101"),
         ("0101010101010110", '0', "011010101010101", "0101010101010101"),
         ("0101010101010110", '0', "011110101010101", "0101010101010101"),
         ("0101010101010101", '1', "001110101010101", "0101010101010110"),
         ("0101010101010101", '1', "001110101010101", "0101010101010101"),
         ("0101010101010110", '1', "010010101010101", "0101010101010101"),
         ("0101010101010110", '1', "010010101010101", "0101010101010110"),
         ("0101010101010110", '0', "000010101010101", "0101010101010101"),
         ("0101010101010110", '0', "000010101010101", "0101010101010101"),
         ("0101010101010110", '0', "000110101010101", "0101010101010101"),
         ("0101010101010110", '0', "001010101010101", "0101010101010101"),
         ("0101010101010110", '0', "001110101010101", "0101010101010101"),
         ("0101010101010110", '0', "010010101010101", "0101010101010110"),
         ("0101010101010110", '0', "010110101010101", "0101010101010101"),
         ("0101010101010110", '0', "011010101010101", "0101010101010101"),
         ("0101010101010110", '0', "011110101010101", "0101010101010101"),
         ("0101010101010101", '1', "010010101010101", "0101010101010110"),
         ("0101010101010101", '1', "010010101010101", "0101010101010101"),
         ("0101010101010110", '1', "010110101010101", "0101010101010101"),
         ("0101010101010110", '1', "010110101010101", "0101010101010110"),
         ("0101010101010110", '0', "000010101010101", "0101010101010101"),
         ("0101010101010110", '0', "000010101010101", "0101010101010101"),
         ("0101010101010110", '0', "000110101010101", "0101010101010101"),
         ("0101010101010110", '0', "001010101010101", "0101010101010101"),
         ("0101010101010110", '0', "001110101010101", "0101010101010101"),
         ("0101010101010110", '0', "010010101010101", "0101010101010101"),
         ("0101010101010110", '0', "010110101010101", "0101010101010110"),
         ("0101010101010110", '0', "011010101010101", "0101010101010101"),
         ("0101010101010110", '0', "011110101010101", "0101010101010101"),
         ("0101010101010101", '1', "010110101010101", "0101010101010110"),
         ("0101010101010101", '1', "010110101010101", "0101010101010101"),
         ("0101010101010110", '1', "011010101010101", "0101010101010101"),
         ("0101010101010110", '1', "011010101010101", "0101010101010110"),
         ("0101010101010110", '0', "000010101010101", "0101010101010101"),
         ("0101010101010110", '0', "000010101010101", "0101010101010101"),
         ("0101010101010110", '0', "000110101010101", "0101010101010101"),
         ("0101010101010110", '0', "001010101010101", "0101010101010101"),
         ("0101010101010110", '0', "001110101010101", "0101010101010101"),
         ("0101010101010110", '0', "010010101010101", "0101010101010101"),
         ("0101010101010110", '0', "010110101010101", "0101010101010101"),
         ("0101010101010110", '0', "011010101010101", "0101010101010110"),
         ("0101010101010110", '0', "011110101010101", "0101010101010101"),
         ("0101010101010101", '1', "011010101010101", "0101010101010110"),
         ("0101010101010101", '1', "011010101010101", "0101010101010101"),
         ("0101010101010110", '1', "011110101010101", "0101010101010101"),
         ("0101010101010110", '1', "011110101010101", "0101010101010110"),
         ("0101010101010110", '0', "000010101010101", "0101010101010101"),
         ("0101010101010110", '0', "000010101010101", "0101010101010101"),
         ("0101010101010110", '0', "000110101010101", "0101010101010101"),
         ("0101010101010110", '0', "001010101010101", "0101010101010101"),
         ("0101010101010110", '0', "001110101010101", "0101010101010101"),
         ("0101010101010110", '0', "010010101010101", "0101010101010101"),
         ("0101010101010110", '0', "010110101010101", "0101010101010101"),
         ("0101010101010110", '0', "011010101010101", "0101010101010101"),
         ("0101010101010110", '0', "011110101010101", "0101010101010110"),
         ("0101010101010101", '1', "011110101010101", "0101010101010110"),
         ("0101010101010101", '1', "011110101010101", "0101010101010101"),
         ("0101010101010101", '0', "000010101010101", "0101010101010101"),
         ("0101010101010101", '0', "000010101010101", "0101010101010101"),
         ("0101010101010101", '0', "000110101010101", "0101010101010101"),
         ("0101010101010101", '0', "001010101010101", "0101010101010101"),
         ("0101010101010101", '0', "001110101010101", "0101010101010101"),
         ("0101010101010101", '0', "010010101010101", "0101010101010101"),
         ("0101010101010101", '0', "010110101010101", "0101010101010101"),
         ("0101010101010101", '0', "011010101010101", "0101010101010101"),
         ("0101010101010101", '0', "011110101010101", "0101010101010101"));
         
   begin
      --  Check each pattern.
      for i in patterns'range loop
         --  Set the inputs.
        d <= patterns(i).d;
        load <= patterns(i).load;
        address <= patterns(i).address;
        wait for 0.25 ns;
        --  Check the outputs.
        assert cout = patterns(i).cout
          report "bad data, memory problem" severity error;
        wait for 0.75 ns;
     end loop;
     -- End the clock
     finish <= '1';
     assert false report "end of test" severity note;
     --  Wait forever; this will finish the simulation.
     wait;
  end process;
end ram16k_tb_arch;
