-- (C) Copyright Collin J. Doering 2015
--
-- This program is free software: you can redistribute it and/or modify
-- it under the terms of the GNU General Public License as published by
-- the Free Software Foundation, either version 3 of the License, or
-- (at your option) any later version.
--
-- This program is distributed in the hope that it will be useful,
-- but WITHOUT ANY WARRANTY; without even the implied warranty of
-- MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
-- GNU General Public License for more details.
--
-- You should have received a copy of the GNU General Public License
-- along with this program.  If not, see <http://www.gnu.org/licenses/>.

-- File: dbit.vhdl
-- Author: Collin J. Doering <collin.doering@rekahsoft.ca>
-- Date: May 22, 2015

library IEEE;
use IEEE.std_logic_1164.all;

entity dbit is
  port (d, load, clk : in  std_logic;
        cout         : out std_logic);
end dbit;

architecture dbit_arch of dbit is
  component mux
    port (a, b, sel : in  std_logic;
          cout      : out std_logic);
  end component;
  component dff
    port (d, clk : in  std_logic;
          cout   : out std_logic);
  end component;

  signal dffOut, muxOut : std_logic;
begin
  MUX_0: mux port map (dffOut, d, load, muxOut);
  DFF_0: dff port map (muxOut, clk, dffOut);
  cout <= dffOut;
end dbit_arch;
