-- (C) Copyright Collin J. Doering 2015
--
-- This program is free software: you can redistribute it and/or modify
-- it under the terms of the GNU General Public License as published by
-- the Free Software Foundation, either version 3 of the License, or
-- (at your option) any later version.
--
-- This program is distributed in the hope that it will be useful,
-- but WITHOUT ANY WARRANTY; without even the implied warranty of
-- MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
-- GNU General Public License for more details.
--
-- You should have received a copy of the GNU General Public License
-- along with this program.  If not, see <http://www.gnu.org/licenses/>.

-- File: ram512_tb.vhdl
-- Author: Collin J. Doering <collin.doering@rekahsoft.ca>
-- Date: May 22, 2015

library IEEE;
use IEEE.std_logic_1164.all;

--  A testbench has no ports.
entity ram512_tb is
end ram512_tb;

architecture ram512_tb_arch of ram512_tb is
   --  Declaration of the component that will be instantiated.
   component ram512
     port (d       : in  std_logic_vector(15 downto 0);
           load    : in  std_logic;
           address : in  std_logic_vector(8 downto 0);
           clk     : in  std_logic;
           cout    : out std_logic_vector(15 downto 0));
   end component;

   -- Declaration of the clock
   component Clock
     port (finish : in  std_logic;
           cout   : out std_logic);
   end component;

   --  Specifies which entity is bound with the component.
   for ram512_0: ram512 use entity work.ram512;

   -- Signals
   signal d, cout           : std_logic_vector(15 downto 0);
   signal address           : std_logic_vector(8 downto 0);
   signal load, finish, clk : std_logic;
begin
  --  Component instantiation.
  OSC_CLK: Clock port map (finish, clk);
  ram512_0: ram512 port map (d, load, address, clk, cout);

   --  This process does the real job.
   process
      type pattern_type is record
         --  The inputs of the ram512.
        d       : std_logic_vector(15 downto 0);
        load    : std_logic;
        address : std_logic_vector(8 downto 0);
        --  The output of the ram512.
        cout    : std_logic_vector(15 downto 0);
      end record;
      --  The patterns to apply.
      type pattern_array is array (natural range <>) of pattern_type;
      constant patterns : pattern_array :=
        (("0000000000000000", '0', "000000000", "0000000000000000"),
         ("0000000000000000", '0', "000000000", "0000000000000000"),
         ("0000000000000000", '1', "000000000", "0000000000000000"),
         ("0000000000000000", '1', "000000000", "0000000000000000"),
         ("0011001100101011", '0', "000000000", "0000000000000000"),
         ("0011001100101011", '0', "000000000", "0000000000000000"),
         ("0011001100101011", '1', "010000010", "0000000000000000"),
         ("0011001100101011", '1', "010000010", "0011001100101011"),
         ("0011001100101011", '0', "000000000", "0000000000000000"),
         ("0011001100101011", '0', "000000000", "0000000000000000"),
         ("0001001001111001", '0', "111011000", "0000000000000000"),
         ("0001001001111001", '0', "111011000", "0000000000000000"),
         ("0001001001111001", '1', "111011000", "0000000000000000"),
         ("0001001001111001", '1', "111011000", "0001001001111001"),
         ("0001001001111001", '0', "111011000", "0001001001111001"),
         ("0001001001111001", '0', "111011000", "0001001001111001"),
         ("0001001001111001", '0', "010000010", "0011001100101011"),
         ("0001001111111111", '0', "010000010", "0011001100101011"),
         ("0001001111111111", '0', "010000010", "0011001100101011"),
         ("0001001111111111", '1', "111111111", "0000000000000000"),
         ("0001001111111111", '1', "111111111", "0001001111111111"),
         ("0001001111111111", '0', "111111111", "0001001111111111"),
         ("0001001111111111", '0', "111111111", "0001001111111111"),
         ("0001001111111111", '0', "111011000", "0001001001111001"),
         ("0001001111111111", '0', "111111111", "0001001111111111"),
         ("0001001111111111", '0', "010101000", "0000000000000000"),
         ("0001001111111111", '0', "010101000", "0000000000000000"),
         ("0001001111111111", '0', "010101001", "0000000000000000"),
         ("0001001111111111", '0', "010101010", "0000000000000000"),
         ("0001001111111111", '0', "010101011", "0000000000000000"),
         ("0001001111111111", '0', "010101100", "0000000000000000"),
         ("0001001111111111", '0', "010101101", "0000000000000000"),
         ("0001001111111111", '0', "010101110", "0000000000000000"),
         ("0001001111111111", '0', "010101111", "0000000000000000"),
         ("0101010101010101", '1', "010101000", "0000000000000000"),
         ("0101010101010101", '1', "010101000", "0101010101010101"),
         ("0101010101010101", '1', "010101001", "0000000000000000"),
         ("0101010101010101", '1', "010101001", "0101010101010101"),
         ("0101010101010101", '1', "010101010", "0000000000000000"),
         ("0101010101010101", '1', "010101010", "0101010101010101"),
         ("0101010101010101", '1', "010101011", "0000000000000000"),
         ("0101010101010101", '1', "010101011", "0101010101010101"),
         ("0101010101010101", '1', "010101100", "0000000000000000"),
         ("0101010101010101", '1', "010101100", "0101010101010101"),
         ("0101010101010101", '1', "010101101", "0000000000000000"),
         ("0101010101010101", '1', "010101101", "0101010101010101"),
         ("0101010101010101", '1', "010101110", "0000000000000000"),
         ("0101010101010101", '1', "010101110", "0101010101010101"),
         ("0101010101010101", '1', "010101111", "0000000000000000"),
         ("0101010101010101", '1', "010101111", "0101010101010101"),
         ("0101010101010101", '0', "010101000", "0101010101010101"),
         ("0101010101010101", '0', "010101000", "0101010101010101"),
         ("0101010101010101", '0', "010101001", "0101010101010101"),
         ("0101010101010101", '0', "010101010", "0101010101010101"),
         ("0101010101010101", '0', "010101011", "0101010101010101"),
         ("0101010101010101", '0', "010101100", "0101010101010101"),
         ("0101010101010101", '0', "010101101", "0101010101010101"),
         ("0101010101010101", '0', "010101110", "0101010101010101"),
         ("0101010101010101", '0', "010101111", "0101010101010101"),
         ("0101010101010110", '1', "010101000", "0101010101010101"),
         ("0101010101010110", '1', "010101000", "0101010101010110"),
         ("0101010101010110", '0', "010101000", "0101010101010110"),
         ("0101010101010110", '0', "010101000", "0101010101010110"),
         ("0101010101010110", '0', "010101001", "0101010101010101"),
         ("0101010101010110", '0', "010101010", "0101010101010101"),
         ("0101010101010110", '0', "010101011", "0101010101010101"),
         ("0101010101010110", '0', "010101100", "0101010101010101"),
         ("0101010101010110", '0', "010101101", "0101010101010101"),
         ("0101010101010110", '0', "010101110", "0101010101010101"),
         ("0101010101010110", '0', "010101111", "0101010101010101"),
         ("0101010101010101", '1', "010101000", "0101010101010110"),
         ("0101010101010101", '1', "010101000", "0101010101010101"),
         ("0101010101010110", '1', "010101001", "0101010101010101"),
         ("0101010101010110", '1', "010101001", "0101010101010110"),
         ("0101010101010110", '0', "010101000", "0101010101010101"),
         ("0101010101010110", '0', "010101000", "0101010101010101"),
         ("0101010101010110", '0', "010101001", "0101010101010110"),
         ("0101010101010110", '0', "010101010", "0101010101010101"),
         ("0101010101010110", '0', "010101011", "0101010101010101"),
         ("0101010101010110", '0', "010101100", "0101010101010101"),
         ("0101010101010110", '0', "010101101", "0101010101010101"),
         ("0101010101010110", '0', "010101110", "0101010101010101"),
         ("0101010101010110", '0', "010101111", "0101010101010101"),
         ("0101010101010101", '1', "010101001", "0101010101010110"),
         ("0101010101010101", '1', "010101001", "0101010101010101"),
         ("0101010101010110", '1', "010101010", "0101010101010101"),
         ("0101010101010110", '1', "010101010", "0101010101010110"),
         ("0101010101010110", '0', "010101000", "0101010101010101"),
         ("0101010101010110", '0', "010101000", "0101010101010101"),
         ("0101010101010110", '0', "010101001", "0101010101010101"),
         ("0101010101010110", '0', "010101010", "0101010101010110"),
         ("0101010101010110", '0', "010101011", "0101010101010101"),
         ("0101010101010110", '0', "010101100", "0101010101010101"),
         ("0101010101010110", '0', "010101101", "0101010101010101"),
         ("0101010101010110", '0', "010101110", "0101010101010101"),
         ("0101010101010110", '0', "010101111", "0101010101010101"),
         ("0101010101010101", '1', "010101010", "0101010101010110"),
         ("0101010101010101", '1', "010101010", "0101010101010101"),
         ("0101010101010110", '1', "010101011", "0101010101010101"),
         ("0101010101010110", '1', "010101011", "0101010101010110"),
         ("0101010101010110", '0', "010101000", "0101010101010101"),
         ("0101010101010110", '0', "010101000", "0101010101010101"),
         ("0101010101010110", '0', "010101001", "0101010101010101"),
         ("0101010101010110", '0', "010101010", "0101010101010101"),
         ("0101010101010110", '0', "010101011", "0101010101010110"),
         ("0101010101010110", '0', "010101100", "0101010101010101"),
         ("0101010101010110", '0', "010101101", "0101010101010101"),
         ("0101010101010110", '0', "010101110", "0101010101010101"),
         ("0101010101010110", '0', "010101111", "0101010101010101"),
         ("0101010101010101", '1', "010101011", "0101010101010110"),
         ("0101010101010101", '1', "010101011", "0101010101010101"),
         ("0101010101010110", '1', "010101100", "0101010101010101"),
         ("0101010101010110", '1', "010101100", "0101010101010110"),
         ("0101010101010110", '0', "010101000", "0101010101010101"),
         ("0101010101010110", '0', "010101000", "0101010101010101"),
         ("0101010101010110", '0', "010101001", "0101010101010101"),
         ("0101010101010110", '0', "010101010", "0101010101010101"),
         ("0101010101010110", '0', "010101011", "0101010101010101"),
         ("0101010101010110", '0', "010101100", "0101010101010110"),
         ("0101010101010110", '0', "010101101", "0101010101010101"),
         ("0101010101010110", '0', "010101110", "0101010101010101"),
         ("0101010101010110", '0', "010101111", "0101010101010101"),
         ("0101010101010101", '1', "010101100", "0101010101010110"),
         ("0101010101010101", '1', "010101100", "0101010101010101"),
         ("0101010101010110", '1', "010101101", "0101010101010101"),
         ("0101010101010110", '1', "010101101", "0101010101010110"),
         ("0101010101010110", '0', "010101000", "0101010101010101"),
         ("0101010101010110", '0', "010101000", "0101010101010101"),
         ("0101010101010110", '0', "010101001", "0101010101010101"),
         ("0101010101010110", '0', "010101010", "0101010101010101"),
         ("0101010101010110", '0', "010101011", "0101010101010101"),
         ("0101010101010110", '0', "010101100", "0101010101010101"),
         ("0101010101010110", '0', "010101101", "0101010101010110"),
         ("0101010101010110", '0', "010101110", "0101010101010101"),
         ("0101010101010110", '0', "010101111", "0101010101010101"),
         ("0101010101010101", '1', "010101101", "0101010101010110"),
         ("0101010101010101", '1', "010101101", "0101010101010101"),
         ("0101010101010110", '1', "010101110", "0101010101010101"),
         ("0101010101010110", '1', "010101110", "0101010101010110"),
         ("0101010101010110", '0', "010101000", "0101010101010101"),
         ("0101010101010110", '0', "010101000", "0101010101010101"),
         ("0101010101010110", '0', "010101001", "0101010101010101"),
         ("0101010101010110", '0', "010101010", "0101010101010101"),
         ("0101010101010110", '0', "010101011", "0101010101010101"),
         ("0101010101010110", '0', "010101100", "0101010101010101"),
         ("0101010101010110", '0', "010101101", "0101010101010101"),
         ("0101010101010110", '0', "010101110", "0101010101010110"),
         ("0101010101010110", '0', "010101111", "0101010101010101"),
         ("0101010101010101", '1', "010101110", "0101010101010110"),
         ("0101010101010101", '1', "010101110", "0101010101010101"),
         ("0101010101010110", '1', "010101111", "0101010101010101"),
         ("0101010101010110", '1', "010101111", "0101010101010110"),
         ("0101010101010110", '0', "010101000", "0101010101010101"),
         ("0101010101010110", '0', "010101000", "0101010101010101"),
         ("0101010101010110", '0', "010101001", "0101010101010101"),
         ("0101010101010110", '0', "010101010", "0101010101010101"),
         ("0101010101010110", '0', "010101011", "0101010101010101"),
         ("0101010101010110", '0', "010101100", "0101010101010101"),
         ("0101010101010110", '0', "010101101", "0101010101010101"),
         ("0101010101010110", '0', "010101110", "0101010101010101"),
         ("0101010101010110", '0', "010101111", "0101010101010110"),
         ("0101010101010101", '1', "010101111", "0101010101010110"),
         ("0101010101010101", '1', "010101111", "0101010101010101"),
         ("0101010101010101", '0', "010101000", "0101010101010101"),
         ("0101010101010101", '0', "010101000", "0101010101010101"),
         ("0101010101010101", '0', "010101001", "0101010101010101"),
         ("0101010101010101", '0', "010101010", "0101010101010101"),
         ("0101010101010101", '0', "010101011", "0101010101010101"),
         ("0101010101010101", '0', "010101100", "0101010101010101"),
         ("0101010101010101", '0', "010101101", "0101010101010101"),
         ("0101010101010101", '0', "010101110", "0101010101010101"),
         ("0101010101010101", '0', "010101111", "0101010101010101"),
         ("0101010101010101", '0', "000101010", "0000000000000000"),
         ("0101010101010101", '0', "000101010", "0000000000000000"),
         ("0101010101010101", '0', "001101010", "0000000000000000"),
         ("0101010101010101", '0', "010101010", "0101010101010101"),
         ("0101010101010101", '0', "011101010", "0000000000000000"),
         ("0101010101010101", '0', "100101010", "0000000000000000"),
         ("0101010101010101", '0', "101101010", "0000000000000000"),
         ("0101010101010101", '0', "110101010", "0000000000000000"),
         ("0101010101010101", '0', "111101010", "0000000000000000"),
         ("0101010101010101", '1', "000101010", "0000000000000000"),
         ("0101010101010101", '1', "000101010", "0101010101010101"),
         ("0101010101010101", '1', "001101010", "0000000000000000"),
         ("0101010101010101", '1', "001101010", "0101010101010101"),
         ("0101010101010101", '1', "010101010", "0101010101010101"),
         ("0101010101010101", '1', "010101010", "0101010101010101"),
         ("0101010101010101", '1', "011101010", "0000000000000000"),
         ("0101010101010101", '1', "011101010", "0101010101010101"),
         ("0101010101010101", '1', "100101010", "0000000000000000"),
         ("0101010101010101", '1', "100101010", "0101010101010101"),
         ("0101010101010101", '1', "101101010", "0000000000000000"),
         ("0101010101010101", '1', "101101010", "0101010101010101"),
         ("0101010101010101", '1', "110101010", "0000000000000000"),
         ("0101010101010101", '1', "110101010", "0101010101010101"),
         ("0101010101010101", '1', "111101010", "0000000000000000"),
         ("0101010101010101", '1', "111101010", "0101010101010101"),
         ("0101010101010101", '0', "000101010", "0101010101010101"),
         ("0101010101010101", '0', "000101010", "0101010101010101"),
         ("0101010101010101", '0', "001101010", "0101010101010101"),
         ("0101010101010101", '0', "010101010", "0101010101010101"),
         ("0101010101010101", '0', "011101010", "0101010101010101"),
         ("0101010101010101", '0', "100101010", "0101010101010101"),
         ("0101010101010101", '0', "101101010", "0101010101010101"),
         ("0101010101010101", '0', "110101010", "0101010101010101"),
         ("0101010101010101", '0', "111101010", "0101010101010101"),
         ("0101010101010110", '1', "000101010", "0101010101010101"),
         ("0101010101010110", '1', "000101010", "0101010101010110"),
         ("0101010101010110", '0', "000101010", "0101010101010110"),
         ("0101010101010110", '0', "000101010", "0101010101010110"),
         ("0101010101010110", '0', "001101010", "0101010101010101"),
         ("0101010101010110", '0', "010101010", "0101010101010101"),
         ("0101010101010110", '0', "011101010", "0101010101010101"),
         ("0101010101010110", '0', "100101010", "0101010101010101"),
         ("0101010101010110", '0', "101101010", "0101010101010101"),
         ("0101010101010110", '0', "110101010", "0101010101010101"),
         ("0101010101010110", '0', "111101010", "0101010101010101"),
         ("0101010101010101", '1', "000101010", "0101010101010110"),
         ("0101010101010101", '1', "000101010", "0101010101010101"),
         ("0101010101010110", '1', "001101010", "0101010101010101"),
         ("0101010101010110", '1', "001101010", "0101010101010110"),
         ("0101010101010110", '0', "000101010", "0101010101010101"),
         ("0101010101010110", '0', "000101010", "0101010101010101"),
         ("0101010101010110", '0', "001101010", "0101010101010110"),
         ("0101010101010110", '0', "010101010", "0101010101010101"),
         ("0101010101010110", '0', "011101010", "0101010101010101"),
         ("0101010101010110", '0', "100101010", "0101010101010101"),
         ("0101010101010110", '0', "101101010", "0101010101010101"),
         ("0101010101010110", '0', "110101010", "0101010101010101"),
         ("0101010101010110", '0', "111101010", "0101010101010101"),
         ("0101010101010101", '1', "001101010", "0101010101010110"),
         ("0101010101010101", '1', "001101010", "0101010101010101"),
         ("0101010101010110", '1', "010101010", "0101010101010101"),
         ("0101010101010110", '1', "010101010", "0101010101010110"),
         ("0101010101010110", '0', "000101010", "0101010101010101"),
         ("0101010101010110", '0', "000101010", "0101010101010101"),
         ("0101010101010110", '0', "001101010", "0101010101010101"),
         ("0101010101010110", '0', "010101010", "0101010101010110"),
         ("0101010101010110", '0', "011101010", "0101010101010101"),
         ("0101010101010110", '0', "100101010", "0101010101010101"),
         ("0101010101010110", '0', "101101010", "0101010101010101"),
         ("0101010101010110", '0', "110101010", "0101010101010101"),
         ("0101010101010110", '0', "111101010", "0101010101010101"),
         ("0101010101010101", '1', "010101010", "0101010101010110"),
         ("0101010101010101", '1', "010101010", "0101010101010101"),
         ("0101010101010110", '1', "011101010", "0101010101010101"),
         ("0101010101010110", '1', "011101010", "0101010101010110"),
         ("0101010101010110", '0', "000101010", "0101010101010101"),
         ("0101010101010110", '0', "000101010", "0101010101010101"),
         ("0101010101010110", '0', "001101010", "0101010101010101"),
         ("0101010101010110", '0', "010101010", "0101010101010101"),
         ("0101010101010110", '0', "011101010", "0101010101010110"),
         ("0101010101010110", '0', "100101010", "0101010101010101"),
         ("0101010101010110", '0', "101101010", "0101010101010101"),
         ("0101010101010110", '0', "110101010", "0101010101010101"),
         ("0101010101010110", '0', "111101010", "0101010101010101"),
         ("0101010101010101", '1', "011101010", "0101010101010110"),
         ("0101010101010101", '1', "011101010", "0101010101010101"),
         ("0101010101010110", '1', "100101010", "0101010101010101"),
         ("0101010101010110", '1', "100101010", "0101010101010110"),
         ("0101010101010110", '0', "000101010", "0101010101010101"),
         ("0101010101010110", '0', "000101010", "0101010101010101"),
         ("0101010101010110", '0', "001101010", "0101010101010101"),
         ("0101010101010110", '0', "010101010", "0101010101010101"),
         ("0101010101010110", '0', "011101010", "0101010101010101"),
         ("0101010101010110", '0', "100101010", "0101010101010110"),
         ("0101010101010110", '0', "101101010", "0101010101010101"),
         ("0101010101010110", '0', "110101010", "0101010101010101"),
         ("0101010101010110", '0', "111101010", "0101010101010101"),
         ("0101010101010101", '1', "100101010", "0101010101010110"),
         ("0101010101010101", '1', "100101010", "0101010101010101"),
         ("0101010101010110", '1', "101101010", "0101010101010101"),
         ("0101010101010110", '1', "101101010", "0101010101010110"),
         ("0101010101010110", '0', "000101010", "0101010101010101"),
         ("0101010101010110", '0', "000101010", "0101010101010101"),
         ("0101010101010110", '0', "001101010", "0101010101010101"),
         ("0101010101010110", '0', "010101010", "0101010101010101"),
         ("0101010101010110", '0', "011101010", "0101010101010101"),
         ("0101010101010110", '0', "100101010", "0101010101010101"),
         ("0101010101010110", '0', "101101010", "0101010101010110"),
         ("0101010101010110", '0', "110101010", "0101010101010101"),
         ("0101010101010110", '0', "111101010", "0101010101010101"),
         ("0101010101010101", '1', "101101010", "0101010101010110"),
         ("0101010101010101", '1', "101101010", "0101010101010101"),
         ("0101010101010110", '1', "110101010", "0101010101010101"),
         ("0101010101010110", '1', "110101010", "0101010101010110"),
         ("0101010101010110", '0', "000101010", "0101010101010101"),
         ("0101010101010110", '0', "000101010", "0101010101010101"),
         ("0101010101010110", '0', "001101010", "0101010101010101"),
         ("0101010101010110", '0', "010101010", "0101010101010101"),
         ("0101010101010110", '0', "011101010", "0101010101010101"),
         ("0101010101010110", '0', "100101010", "0101010101010101"),
         ("0101010101010110", '0', "101101010", "0101010101010101"),
         ("0101010101010110", '0', "110101010", "0101010101010110"),
         ("0101010101010110", '0', "111101010", "0101010101010101"),
         ("0101010101010101", '1', "110101010", "0101010101010110"),
         ("0101010101010101", '1', "110101010", "0101010101010101"),
         ("0101010101010110", '1', "111101010", "0101010101010101"),
         ("0101010101010110", '1', "111101010", "0101010101010110"),
         ("0101010101010110", '0', "000101010", "0101010101010101"),
         ("0101010101010110", '0', "000101010", "0101010101010101"),
         ("0101010101010110", '0', "001101010", "0101010101010101"),
         ("0101010101010110", '0', "010101010", "0101010101010101"),
         ("0101010101010110", '0', "011101010", "0101010101010101"),
         ("0101010101010110", '0', "100101010", "0101010101010101"),
         ("0101010101010110", '0', "101101010", "0101010101010101"),
         ("0101010101010110", '0', "110101010", "0101010101010101"),
         ("0101010101010110", '0', "111101010", "0101010101010110"),
         ("0101010101010101", '1', "111101010", "0101010101010110"),
         ("0101010101010101", '1', "111101010", "0101010101010101"),
         ("0101010101010101", '0', "000101010", "0101010101010101"),
         ("0101010101010101", '0', "000101010", "0101010101010101"),
         ("0101010101010101", '0', "001101010", "0101010101010101"),
         ("0101010101010101", '0', "010101010", "0101010101010101"),
         ("0101010101010101", '0', "011101010", "0101010101010101"),
         ("0101010101010101", '0', "100101010", "0101010101010101"),
         ("0101010101010101", '0', "101101010", "0101010101010101"),
         ("0101010101010101", '0', "110101010", "0101010101010101"),
         ("0101010101010101", '0', "111101010", "0101010101010101"));
         
   begin
      --  Check each pattern.
      for i in patterns'range loop
         --  Set the inputs.
        d <= patterns(i).d;
        load <= patterns(i).load;
        address <= patterns(i).address;
        wait for 0.25 ns;
        --  Check the outputs.
        assert cout = patterns(i).cout
          report "bad data, memory problem" severity error;
        wait for 0.75 ns;
     end loop;
     -- End the clock
     finish <= '1';
     assert false report "end of test" severity note;
     --  Wait forever; this will finish the simulation.
     wait;
  end process;
end ram512_tb_arch;
