library IEEE;
use IEEE.std_logic_1164.all;

--  A testbench has no ports.
entity ram4k_tb is
end ram4k_tb;

architecture ram4k_tb_arch of ram4k_tb is
   --  Declaration of the component that will be instantiated.
   component ram4k
     port (d       : in std_logic_vector(15 downto 0);
           load    : in std_logic;
           address : in std_logic_vector(11 downto 0);
           clk     : in std_logic;
           cout    : out std_logic_vector(15 downto 0));
   end component;
   -- Declaration of the clock
   component Clock
     port (finish : in std_logic;
           cout   : out std_logic);
   end component;
   
   --  Specifies which entity is bound with the component.
   for ram4k_0: ram4k use entity work.ram4k;
   signal d, cout : std_logic_vector(15 downto 0);
   signal address : std_logic_vector(11 downto 0);
   signal load, finish, clk : std_logic;
begin
  --  Component instantiation.
  OSC_CLK: Clock port map (finish, clk);
  ram4k_0: ram4k port map (d, load, address, clk, cout);

   --  This process does the real job.
   process
      type pattern_type is record
         --  The inputs of the ram4k.
        d       : std_logic_vector(15 downto 0);
        load    : std_logic;
        address : std_logic_vector(11 downto 0);
        --  The output of the ram4k.
        cout    : std_logic_vector(15 downto 0);
      end record;
      --  The patterns to apply.
      type pattern_array is array (natural range <>) of pattern_type;
      constant patterns : pattern_array :=
        (("0000000000000000", '0', "000000000000", "0000000000000000"),
         ("0000000000000000", '0', "000000000000", "0000000000000000"),
         ("0000000000000000", '1', "000000000000", "0000000000000000"),
         ("0000000000000000", '1', "000000000000", "0000000000000000"),
         ("0000010001010111", '0', "000000000000", "0000000000000000"),
         ("0000010001010111", '0', "000000000000", "0000000000000000"),
         ("0000010001010111", '1', "010001010111", "0000000000000000"),
         ("0000010001010111", '1', "010001010111", "0000010001010111"),
         ("0000010001010111", '0', "000000000000", "0000000000000000"),
         ("0000010001010111", '0', "000000000000", "0000000000000000"),
         ("0000110110111001", '0', "110110111001", "0000000000000000"),
         ("0000110110111001", '0', "110110111001", "0000000000000000"),
         ("0000110110111001", '1', "110110111001", "0000000000000000"),
         ("0000110110111001", '1', "110110111001", "0000110110111001"),
         ("0000110110111001", '0', "110110111001", "0000110110111001"),
         ("0000110110111001", '0', "110110111001", "0000110110111001"),
         ("0000110110111001", '0', "010001010111", "0000010001010111"),
         ("0000111111111111", '0', "010001010111", "0000010001010111"),
         ("0000111111111111", '0', "010001010111", "0000010001010111"),
         ("0000111111111111", '1', "111111111111", "0000000000000000"),
         ("0000111111111111", '1', "111111111111", "0000111111111111"),
         ("0000111111111111", '0', "111111111111", "0000111111111111"),
         ("0000111111111111", '0', "111111111111", "0000111111111111"),
         ("0000111111111111", '0', "110110111001", "0000110110111001"),
         ("0000111111111111", '0', "111111111111", "0000111111111111"),
         ("0000111111111111", '0', "101010101000", "0000000000000000"),
         ("0000111111111111", '0', "101010101000", "0000000000000000"),
         ("0000111111111111", '0', "101010101001", "0000000000000000"),
         ("0000111111111111", '0', "101010101010", "0000000000000000"),
         ("0000111111111111", '0', "101010101011", "0000000000000000"),
         ("0000111111111111", '0', "101010101100", "0000000000000000"),
         ("0000111111111111", '0', "101010101101", "0000000000000000"),
         ("0000111111111111", '0', "101010101110", "0000000000000000"),
         ("0000111111111111", '0', "101010101111", "0000000000000000"),
         ("0101010101010101", '1', "101010101000", "0000000000000000"),
         ("0101010101010101", '1', "101010101000", "0101010101010101"),
         ("0101010101010101", '1', "101010101001", "0000000000000000"),
         ("0101010101010101", '1', "101010101001", "0101010101010101"),
         ("0101010101010101", '1', "101010101010", "0000000000000000"),
         ("0101010101010101", '1', "101010101010", "0101010101010101"),
         ("0101010101010101", '1', "101010101011", "0000000000000000"),
         ("0101010101010101", '1', "101010101011", "0101010101010101"),
         ("0101010101010101", '1', "101010101100", "0000000000000000"),
         ("0101010101010101", '1', "101010101100", "0101010101010101"),
         ("0101010101010101", '1', "101010101101", "0000000000000000"),
         ("0101010101010101", '1', "101010101101", "0101010101010101"),
         ("0101010101010101", '1', "101010101110", "0000000000000000"),
         ("0101010101010101", '1', "101010101110", "0101010101010101"),
         ("0101010101010101", '1', "101010101111", "0000000000000000"),
         ("0101010101010101", '1', "101010101111", "0101010101010101"),
         ("0101010101010101", '0', "101010101000", "0101010101010101"),
         ("0101010101010101", '0', "101010101000", "0101010101010101"),
         ("0101010101010101", '0', "101010101001", "0101010101010101"),
         ("0101010101010101", '0', "101010101010", "0101010101010101"),
         ("0101010101010101", '0', "101010101011", "0101010101010101"),
         ("0101010101010101", '0', "101010101100", "0101010101010101"),
         ("0101010101010101", '0', "101010101101", "0101010101010101"),
         ("0101010101010101", '0', "101010101110", "0101010101010101"),
         ("0101010101010101", '0', "101010101111", "0101010101010101"),
         ("0101010101010110", '1', "101010101000", "0101010101010101"),
         ("0101010101010110", '1', "101010101000", "0101010101010110"),
         ("0101010101010110", '0', "101010101000", "0101010101010110"),
         ("0101010101010110", '0', "101010101000", "0101010101010110"),
         ("0101010101010110", '0', "101010101001", "0101010101010101"),
         ("0101010101010110", '0', "101010101010", "0101010101010101"),
         ("0101010101010110", '0', "101010101011", "0101010101010101"),
         ("0101010101010110", '0', "101010101100", "0101010101010101"),
         ("0101010101010110", '0', "101010101101", "0101010101010101"),
         ("0101010101010110", '0', "101010101110", "0101010101010101"),
         ("0101010101010110", '0', "101010101111", "0101010101010101"),
         ("0101010101010101", '1', "101010101000", "0101010101010110"),
         ("0101010101010101", '1', "101010101000", "0101010101010101"),
         ("0101010101010110", '1', "101010101001", "0101010101010101"),
         ("0101010101010110", '1', "101010101001", "0101010101010110"),
         ("0101010101010110", '0', "101010101000", "0101010101010101"),
         ("0101010101010110", '0', "101010101000", "0101010101010101"),
         ("0101010101010110", '0', "101010101001", "0101010101010110"),
         ("0101010101010110", '0', "101010101010", "0101010101010101"),
         ("0101010101010110", '0', "101010101011", "0101010101010101"),
         ("0101010101010110", '0', "101010101100", "0101010101010101"),
         ("0101010101010110", '0', "101010101101", "0101010101010101"),
         ("0101010101010110", '0', "101010101110", "0101010101010101"),
         ("0101010101010110", '0', "101010101111", "0101010101010101"),
         ("0101010101010101", '1', "101010101001", "0101010101010110"),
         ("0101010101010101", '1', "101010101001", "0101010101010101"),
         ("0101010101010110", '1', "101010101010", "0101010101010101"),
         ("0101010101010110", '1', "101010101010", "0101010101010110"),
         ("0101010101010110", '0', "101010101000", "0101010101010101"),
         ("0101010101010110", '0', "101010101000", "0101010101010101"),
         ("0101010101010110", '0', "101010101001", "0101010101010101"),
         ("0101010101010110", '0', "101010101010", "0101010101010110"),
         ("0101010101010110", '0', "101010101011", "0101010101010101"),
         ("0101010101010110", '0', "101010101100", "0101010101010101"),
         ("0101010101010110", '0', "101010101101", "0101010101010101"),
         ("0101010101010110", '0', "101010101110", "0101010101010101"),
         ("0101010101010110", '0', "101010101111", "0101010101010101"),
         ("0101010101010101", '1', "101010101010", "0101010101010110"),
         ("0101010101010101", '1', "101010101010", "0101010101010101"),
         ("0101010101010110", '1', "101010101011", "0101010101010101"),
         ("0101010101010110", '1', "101010101011", "0101010101010110"),
         ("0101010101010110", '0', "101010101000", "0101010101010101"),
         ("0101010101010110", '0', "101010101000", "0101010101010101"),
         ("0101010101010110", '0', "101010101001", "0101010101010101"),
         ("0101010101010110", '0', "101010101010", "0101010101010101"),
         ("0101010101010110", '0', "101010101011", "0101010101010110"),
         ("0101010101010110", '0', "101010101100", "0101010101010101"),
         ("0101010101010110", '0', "101010101101", "0101010101010101"),
         ("0101010101010110", '0', "101010101110", "0101010101010101"),
         ("0101010101010110", '0', "101010101111", "0101010101010101"),
         ("0101010101010101", '1', "101010101011", "0101010101010110"),
         ("0101010101010101", '1', "101010101011", "0101010101010101"),
         ("0101010101010110", '1', "101010101100", "0101010101010101"),
         ("0101010101010110", '1', "101010101100", "0101010101010110"),
         ("0101010101010110", '0', "101010101000", "0101010101010101"),
         ("0101010101010110", '0', "101010101000", "0101010101010101"),
         ("0101010101010110", '0', "101010101001", "0101010101010101"),
         ("0101010101010110", '0', "101010101010", "0101010101010101"),
         ("0101010101010110", '0', "101010101011", "0101010101010101"),
         ("0101010101010110", '0', "101010101100", "0101010101010110"),
         ("0101010101010110", '0', "101010101101", "0101010101010101"),
         ("0101010101010110", '0', "101010101110", "0101010101010101"),
         ("0101010101010110", '0', "101010101111", "0101010101010101"),
         ("0101010101010101", '1', "101010101100", "0101010101010110"),
         ("0101010101010101", '1', "101010101100", "0101010101010101"),
         ("0101010101010110", '1', "101010101101", "0101010101010101"),
         ("0101010101010110", '1', "101010101101", "0101010101010110"),
         ("0101010101010110", '0', "101010101000", "0101010101010101"),
         ("0101010101010110", '0', "101010101000", "0101010101010101"),
         ("0101010101010110", '0', "101010101001", "0101010101010101"),
         ("0101010101010110", '0', "101010101010", "0101010101010101"),
         ("0101010101010110", '0', "101010101011", "0101010101010101"),
         ("0101010101010110", '0', "101010101100", "0101010101010101"),
         ("0101010101010110", '0', "101010101101", "0101010101010110"),
         ("0101010101010110", '0', "101010101110", "0101010101010101"),
         ("0101010101010110", '0', "101010101111", "0101010101010101"),
         ("0101010101010101", '1', "101010101101", "0101010101010110"),
         ("0101010101010101", '1', "101010101101", "0101010101010101"),
         ("0101010101010110", '1', "101010101110", "0101010101010101"),
         ("0101010101010110", '1', "101010101110", "0101010101010110"),
         ("0101010101010110", '0', "101010101000", "0101010101010101"),
         ("0101010101010110", '0', "101010101000", "0101010101010101"),
         ("0101010101010110", '0', "101010101001", "0101010101010101"),
         ("0101010101010110", '0', "101010101010", "0101010101010101"),
         ("0101010101010110", '0', "101010101011", "0101010101010101"),
         ("0101010101010110", '0', "101010101100", "0101010101010101"),
         ("0101010101010110", '0', "101010101101", "0101010101010101"),
         ("0101010101010110", '0', "101010101110", "0101010101010110"),
         ("0101010101010110", '0', "101010101111", "0101010101010101"),
         ("0101010101010101", '1', "101010101110", "0101010101010110"),
         ("0101010101010101", '1', "101010101110", "0101010101010101"),
         ("0101010101010110", '1', "101010101111", "0101010101010101"),
         ("0101010101010110", '1', "101010101111", "0101010101010110"),
         ("0101010101010110", '0', "101010101000", "0101010101010101"),
         ("0101010101010110", '0', "101010101000", "0101010101010101"),
         ("0101010101010110", '0', "101010101001", "0101010101010101"),
         ("0101010101010110", '0', "101010101010", "0101010101010101"),
         ("0101010101010110", '0', "101010101011", "0101010101010101"),
         ("0101010101010110", '0', "101010101100", "0101010101010101"),
         ("0101010101010110", '0', "101010101101", "0101010101010101"),
         ("0101010101010110", '0', "101010101110", "0101010101010101"),
         ("0101010101010110", '0', "101010101111", "0101010101010110"),
         ("0101010101010101", '1', "101010101111", "0101010101010110"),
         ("0101010101010101", '1', "101010101111", "0101010101010101"),
         ("0101010101010101", '0', "101010101000", "0101010101010101"),
         ("0101010101010101", '0', "101010101000", "0101010101010101"),
         ("0101010101010101", '0', "101010101001", "0101010101010101"),
         ("0101010101010101", '0', "101010101010", "0101010101010101"),
         ("0101010101010101", '0', "101010101011", "0101010101010101"),
         ("0101010101010101", '0', "101010101100", "0101010101010101"),
         ("0101010101010101", '0', "101010101101", "0101010101010101"),
         ("0101010101010101", '0', "101010101110", "0101010101010101"),
         ("0101010101010101", '0', "101010101111", "0101010101010101"),
         ("0101010101010101", '0', "000101010101", "0000000000000000"),
         ("0101010101010101", '0', "000101010101", "0000000000000000"),
         ("0101010101010101", '0', "001101010101", "0000000000000000"),
         ("0101010101010101", '0', "010101010101", "0000000000000000"),
         ("0101010101010101", '0', "011101010101", "0000000000000000"),
         ("0101010101010101", '0', "100101010101", "0000000000000000"),
         ("0101010101010101", '0', "101101010101", "0000000000000000"),
         ("0101010101010101", '0', "110101010101", "0000000000000000"),
         ("0101010101010101", '0', "111101010101", "0000000000000000"),
         ("0101010101010101", '1', "000101010101", "0000000000000000"),
         ("0101010101010101", '1', "000101010101", "0101010101010101"),
         ("0101010101010101", '1', "001101010101", "0000000000000000"),
         ("0101010101010101", '1', "001101010101", "0101010101010101"),
         ("0101010101010101", '1', "010101010101", "0000000000000000"),
         ("0101010101010101", '1', "010101010101", "0101010101010101"),
         ("0101010101010101", '1', "011101010101", "0000000000000000"),
         ("0101010101010101", '1', "011101010101", "0101010101010101"),
         ("0101010101010101", '1', "100101010101", "0000000000000000"),
         ("0101010101010101", '1', "100101010101", "0101010101010101"),
         ("0101010101010101", '1', "101101010101", "0000000000000000"),
         ("0101010101010101", '1', "101101010101", "0101010101010101"),
         ("0101010101010101", '1', "110101010101", "0000000000000000"),
         ("0101010101010101", '1', "110101010101", "0101010101010101"),
         ("0101010101010101", '1', "111101010101", "0000000000000000"),
         ("0101010101010101", '1', "111101010101", "0101010101010101"),
         ("0101010101010101", '0', "000101010101", "0101010101010101"),
         ("0101010101010101", '0', "000101010101", "0101010101010101"),
         ("0101010101010101", '0', "001101010101", "0101010101010101"),
         ("0101010101010101", '0', "010101010101", "0101010101010101"),
         ("0101010101010101", '0', "011101010101", "0101010101010101"),
         ("0101010101010101", '0', "100101010101", "0101010101010101"),
         ("0101010101010101", '0', "101101010101", "0101010101010101"),
         ("0101010101010101", '0', "110101010101", "0101010101010101"),
         ("0101010101010101", '0', "111101010101", "0101010101010101"),
         ("0101010101010110", '1', "000101010101", "0101010101010101"),
         ("0101010101010110", '1', "000101010101", "0101010101010110"),
         ("0101010101010110", '0', "000101010101", "0101010101010110"),
         ("0101010101010110", '0', "000101010101", "0101010101010110"),
         ("0101010101010110", '0', "001101010101", "0101010101010101"),
         ("0101010101010110", '0', "010101010101", "0101010101010101"),
         ("0101010101010110", '0', "011101010101", "0101010101010101"),
         ("0101010101010110", '0', "100101010101", "0101010101010101"),
         ("0101010101010110", '0', "101101010101", "0101010101010101"),
         ("0101010101010110", '0', "110101010101", "0101010101010101"),
         ("0101010101010110", '0', "111101010101", "0101010101010101"),
         ("0101010101010101", '1', "000101010101", "0101010101010110"),
         ("0101010101010101", '1', "000101010101", "0101010101010101"),
         ("0101010101010110", '1', "001101010101", "0101010101010101"),
         ("0101010101010110", '1', "001101010101", "0101010101010110"),
         ("0101010101010110", '0', "000101010101", "0101010101010101"),
         ("0101010101010110", '0', "000101010101", "0101010101010101"),
         ("0101010101010110", '0', "001101010101", "0101010101010110"),
         ("0101010101010110", '0', "010101010101", "0101010101010101"),
         ("0101010101010110", '0', "011101010101", "0101010101010101"),
         ("0101010101010110", '0', "100101010101", "0101010101010101"),
         ("0101010101010110", '0', "101101010101", "0101010101010101"),
         ("0101010101010110", '0', "110101010101", "0101010101010101"),
         ("0101010101010110", '0', "111101010101", "0101010101010101"),
         ("0101010101010101", '1', "001101010101", "0101010101010110"),
         ("0101010101010101", '1', "001101010101", "0101010101010101"),
         ("0101010101010110", '1', "010101010101", "0101010101010101"),
         ("0101010101010110", '1', "010101010101", "0101010101010110"),
         ("0101010101010110", '0', "000101010101", "0101010101010101"),
         ("0101010101010110", '0', "000101010101", "0101010101010101"),
         ("0101010101010110", '0', "001101010101", "0101010101010101"),
         ("0101010101010110", '0', "010101010101", "0101010101010110"),
         ("0101010101010110", '0', "011101010101", "0101010101010101"),
         ("0101010101010110", '0', "100101010101", "0101010101010101"),
         ("0101010101010110", '0', "101101010101", "0101010101010101"),
         ("0101010101010110", '0', "110101010101", "0101010101010101"),
         ("0101010101010110", '0', "111101010101", "0101010101010101"),
         ("0101010101010101", '1', "010101010101", "0101010101010110"),
         ("0101010101010101", '1', "010101010101", "0101010101010101"),
         ("0101010101010110", '1', "011101010101", "0101010101010101"),
         ("0101010101010110", '1', "011101010101", "0101010101010110"),
         ("0101010101010110", '0', "000101010101", "0101010101010101"),
         ("0101010101010110", '0', "000101010101", "0101010101010101"),
         ("0101010101010110", '0', "001101010101", "0101010101010101"),
         ("0101010101010110", '0', "010101010101", "0101010101010101"),
         ("0101010101010110", '0', "011101010101", "0101010101010110"),
         ("0101010101010110", '0', "100101010101", "0101010101010101"),
         ("0101010101010110", '0', "101101010101", "0101010101010101"),
         ("0101010101010110", '0', "110101010101", "0101010101010101"),
         ("0101010101010110", '0', "111101010101", "0101010101010101"),
         ("0101010101010101", '1', "011101010101", "0101010101010110"),
         ("0101010101010101", '1', "011101010101", "0101010101010101"),
         ("0101010101010110", '1', "100101010101", "0101010101010101"),
         ("0101010101010110", '1', "100101010101", "0101010101010110"),
         ("0101010101010110", '0', "000101010101", "0101010101010101"),
         ("0101010101010110", '0', "000101010101", "0101010101010101"),
         ("0101010101010110", '0', "001101010101", "0101010101010101"),
         ("0101010101010110", '0', "010101010101", "0101010101010101"),
         ("0101010101010110", '0', "011101010101", "0101010101010101"),
         ("0101010101010110", '0', "100101010101", "0101010101010110"),
         ("0101010101010110", '0', "101101010101", "0101010101010101"),
         ("0101010101010110", '0', "110101010101", "0101010101010101"),
         ("0101010101010110", '0', "111101010101", "0101010101010101"),
         ("0101010101010101", '1', "100101010101", "0101010101010110"),
         ("0101010101010101", '1', "100101010101", "0101010101010101"),
         ("0101010101010110", '1', "101101010101", "0101010101010101"),
         ("0101010101010110", '1', "101101010101", "0101010101010110"),
         ("0101010101010110", '0', "000101010101", "0101010101010101"),
         ("0101010101010110", '0', "000101010101", "0101010101010101"),
         ("0101010101010110", '0', "001101010101", "0101010101010101"),
         ("0101010101010110", '0', "010101010101", "0101010101010101"),
         ("0101010101010110", '0', "011101010101", "0101010101010101"),
         ("0101010101010110", '0', "100101010101", "0101010101010101"),
         ("0101010101010110", '0', "101101010101", "0101010101010110"),
         ("0101010101010110", '0', "110101010101", "0101010101010101"),
         ("0101010101010110", '0', "111101010101", "0101010101010101"),
         ("0101010101010101", '1', "101101010101", "0101010101010110"),
         ("0101010101010101", '1', "101101010101", "0101010101010101"),
         ("0101010101010110", '1', "110101010101", "0101010101010101"),
         ("0101010101010110", '1', "110101010101", "0101010101010110"),
         ("0101010101010110", '0', "000101010101", "0101010101010101"),
         ("0101010101010110", '0', "000101010101", "0101010101010101"),
         ("0101010101010110", '0', "001101010101", "0101010101010101"),
         ("0101010101010110", '0', "010101010101", "0101010101010101"),
         ("0101010101010110", '0', "011101010101", "0101010101010101"),
         ("0101010101010110", '0', "100101010101", "0101010101010101"),
         ("0101010101010110", '0', "101101010101", "0101010101010101"),
         ("0101010101010110", '0', "110101010101", "0101010101010110"),
         ("0101010101010110", '0', "111101010101", "0101010101010101"),
         ("0101010101010101", '1', "110101010101", "0101010101010110"),
         ("0101010101010101", '1', "110101010101", "0101010101010101"),
         ("0101010101010110", '1', "111101010101", "0101010101010101"),
         ("0101010101010110", '1', "111101010101", "0101010101010110"),
         ("0101010101010110", '0', "000101010101", "0101010101010101"),
         ("0101010101010110", '0', "000101010101", "0101010101010101"),
         ("0101010101010110", '0', "001101010101", "0101010101010101"),
         ("0101010101010110", '0', "010101010101", "0101010101010101"),
         ("0101010101010110", '0', "011101010101", "0101010101010101"),
         ("0101010101010110", '0', "100101010101", "0101010101010101"),
         ("0101010101010110", '0', "101101010101", "0101010101010101"),
         ("0101010101010110", '0', "110101010101", "0101010101010101"),
         ("0101010101010110", '0', "111101010101", "0101010101010110"),
         ("0101010101010101", '1', "111101010101", "0101010101010110"),
         ("0101010101010101", '1', "111101010101", "0101010101010101"),
         ("0101010101010101", '0', "000101010101", "0101010101010101"),
         ("0101010101010101", '0', "000101010101", "0101010101010101"),
         ("0101010101010101", '0', "001101010101", "0101010101010101"),
         ("0101010101010101", '0', "010101010101", "0101010101010101"),
         ("0101010101010101", '0', "011101010101", "0101010101010101"),
         ("0101010101010101", '0', "100101010101", "0101010101010101"),
         ("0101010101010101", '0', "101101010101", "0101010101010101"),
         ("0101010101010101", '0', "110101010101", "0101010101010101"),
         ("0101010101010101", '0', "111101010101", "0101010101010101"));
         
   begin
      --  Check each pattern.
      for i in patterns'range loop
         --  Set the inputs.
        d <= patterns(i).d;
        load <= patterns(i).load;
        address <= patterns(i).address;
        wait for 0.25 ns;
        --  Check the outputs.
        assert cout = patterns(i).cout
          report "bad data, memory problem" severity error;
        wait for 0.75 ns;
     end loop;
     -- End the clock
     finish <= '1';
     assert false report "end of test" severity note;
     --  Wait forever; this will finish the simulation.
     wait;
  end process;
end ram4k_tb_arch;
