-- (C) Copyright Collin J. Doering 2015
--
-- This program is free software: you can redistribute it and/or modify
-- it under the terms of the GNU General Public License as published by
-- the Free Software Foundation, either version 3 of the License, or
-- (at your option) any later version.
--
-- This program is distributed in the hope that it will be useful,
-- but WITHOUT ANY WARRANTY; without even the implied warranty of
-- MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
-- GNU General Public License for more details.
--
-- You should have received a copy of the GNU General Public License
-- along with this program.  If not, see <http://www.gnu.org/licenses/>.

-- File: cpu_tb.vhdl
-- Author: Collin J. Doering <collin.doering@rekahsoft.ca>
-- Date: May 22, 2015

library IEEE;
use IEEE.std_logic_1164.all;

--  A testbench has no ports.
entity cpu_tb is
end cpu_tb;
architecture cpu_tb_arch of cpu_tb is
   --  Declaration of the component that will be instantiated.
   component cpu
     port (inM, instruction : in  std_logic_vector(15 downto 0);
           reset, clk       : in  std_logic;
           outM             : out std_logic_vector(15 downto 0);
           writeM           : out std_logic;
           addressM, pcOut  : out std_logic_vector(14 downto 0));
   end component;

   -- Declaration of the clock
   component Clock
     port (finish : in  std_logic;
           cout   : out std_logic);
   end component;
   
   --  Specifies which entity is bound with the component.
   for cpu_0: cpu use entity work.cpu;

   -- Signals
   signal reset, writeM, finish, clk : std_logic;
   signal inM, instruction, outM     : std_logic_vector(15 downto 0);
   signal addressM, pcOut            : std_logic_vector(14 downto 0);

   --signal regd : <<signal regDOut : std_logic_vector(15 downto 0)>>;
begin
  --  Component instantiation.
  OSC_CLK: Clock port map (finish, clk);
  cpu_0: cpu port map (inM, instruction, reset, clk, outM, writeM, addressM, pcOut);

   --  This process does the real job.
   process
      type pattern_type is record
         --  The inputs of the cpu.
         inM, instruction : std_logic_vector(15 downto 0);
         reset            : std_logic;
         --  The output of the cpu.
         outM             : std_logic_vector(15 downto 0);
         writeM           : std_logic;
         addressM, pcOut  : std_logic_vector(14 downto 0);
         registerD        : std_logic_vector(15 downto 0);
         -- dregister TODO
      end record;
      --  The patterns to apply.
      type pattern_array is array (natural range <>) of pattern_type;
      -- Below many checks fail, due to syncronization (the compare data given
      -- by the nand to tetris course uses a two phase clock (??) whereas this
      -- implementation uses a single pase. This still needs to be confirmed
      -- and if it is the case, have the test data modified accoridingly.
      constant patterns : pattern_array :=
        (("0000000000000000", "0011000000111001", '0', "----------------", '0', "000000000000000", "000000000000000", "0000000000000000"), -- 0
      -- ("0000"            , "3039"            , '0', "0000"            , '0', "0000"           , "0000"           , "0000"            )
         ("0000000000000000", "0011000000111001", '0', "----------------", '0', "011000000111001", "000000000000001", "0000000000000000"), -- 1
      -- ("0000"            , "3039"            , '0', "0000"            , '0', "3039"           , "0001"           , "0000"            )
         ("0000000000000000", "1110110000010000", '0', "----------------", '0', "011000000111001", "000000000000001", "0011000000111001"), -- 2 (fails: pc)
      -- ("0000"            , "EC10"            , '0', "0000"            , '0', "3039"           , "0001"           , "3039"            )
         ("0000000000000000", "1110110000010000", '0', "----------------", '0', "011000000111001", "000000000000010", "0011000000111001"), -- 3 (fails: pc)
      -- ("0000"            , "EC10"            , '0', "0000"            , '0', "3039"           , "0002"           , "3039"            )
         ("0000000000000000", "0101101110100000", '0', "----------------", '0', "011000000111001", "000000000000010", "0011000000111001"), -- 4 (fails: pc)
      -- ("0000"            , "5BA0"            , '0', "0000"            , '0', "3039"           , "0002"           , "3039"            )
         ("0000000000000000", "0101101110100000", '0', "----------------", '0', "101101110100000", "000000000000011", "0011000000111001"), -- 5 (fails: pc)
      -- ("0000"            , "5BA0"            , '0', "0000"            , '0', "5BA0"           , "0003"           , "3039"            )
         ("0000000000000000", "1110000111010000", '0', "----------------", '0', "101101110100000", "000000000000011", "0010101101100111"), -- 6 (fails: pc)
      -- ("0000"            , "E1D0"            , '0', "0000"            , '0', "5BA0"           , "0003"           , "2B67"            )
         ("0000000000000000", "1110000111010000", '0', "----------------", '0', "101101110100000", "000000000000100", "0010101101100111"), -- 7 (fails: pc)
      -- ("0000"            , "E1D0"            , '0', "0000"            , '0', "5BA0"           , "0004"           , "2B67"            )
         ("0000000000000000", "0000001111101000", '0', "----------------", '0', "101101110100000", "000000000000100", "0010101101100111"), -- 8 (fails: pc)
      -- ("0000"            , "03E8"            , '0', "0000"            , '0', "5BA0"           , "0004"           , "2B67"            )
         ("0000000000000000", "0000001111101000", '0', "----------------", '0', "000001111101000", "000000000000101", "0010101101100111"), -- 9 (fails: pc)
      -- ("0000"            , "03E8"            , '0', "0000"            , '0', "03E8"           , "0005"           , "2B67"            )
         ("0000000000000000", "1110001100001000", '0', "0010101101100111", '1', "000001111101000", "000000000000101", "0010101101100111"), -- 10 (fails: cpu pc)
      -- ("0000"            , "E308"            , '0', "2B67"            , '1', "03E8"           , "0005"           , "2B67"            )
         ("0000000000000000", "1110001100001000", '0', "0010101101100111", '1', "000001111101000", "000000000000110", "0010101101100111"), -- 11 (fails: cpu pc)
      -- ("0000"            , "E308"            , '0', "2B67"            , '1', "03E8"           , "0006"           , "2B67"            )
         ("0000000000000000", "0000001111101001", '0', "----------------", '0', "000001111101000", "000000000000110", "0010101101100111"), -- 12 (fails: pc)
      -- ("0000"            , "03E9"            , '0', "0000"            , '0', "03E8"           , "0006"           , "2B67"            )
         ("0000000000000000", "0000001111101001", '0', "----------------", '0', "000001111101001", "000000000000111", "0010101101100111"), -- 13 (fails: pc)
      -- ("0000"            , "03E9"            , '0', "0000"            , '0', "03E9"           , "0007"           , "2B67"            )
         ("0000000000000000", "1110001110011000", '0', "0010101101100110", '1', "000001111101001", "000000000000111", "0010101101100110"), -- 14 (fails: cpu pc)
      -- ("0000"            , "E398"            , '0', "2B66"            , '1', "03E9"           , "0007"           , "2B66"            )
         ("0000000000000000", "1110001110011000", '0', "0010101101100101", '1', "000001111101001", "000000000001000", "0010101101100110"), -- 15 (fails: cpu pc)
      -- ("0000"            , "E398"            , '0', "2B65"            , '1', "03E9"           , "0008"           , "2B66"            )
         ("0000000000000000", "0000001111101000", '0', "----------------", '0', "000001111101001", "000000000001000", "0010101101100110"), -- 16 (fails: pc)
      -- ("0000"            , "03E8"            , '0', "0000"            , '0', "03E9"           , "0008"           , "2B66"            )
         ("0000000000000000", "0000001111101000", '0', "----------------", '0', "000001111101000", "000000000001001", "0010101101100110"), -- 17 (fails: pc)
      -- ("0000"            , "03E8"            , '0', "0000"            , '0', "03E8"           , "0009"           , "2B66"            )
         ("0010101101100111", "1111010011010000", '0', "----------------", '0', "000001111101000", "000000000001001", "1111111111111111"), -- 18 (fails: pc)
      -- ("2B67"            , "F4D0"            , '0', "0000"            , '0', "03E8"           , "0009"           , "FFFF"            )
         ("0010101101100111", "1111010011010000", '0', "----------------", '0', "000001111101000", "000000000001010", "1111111111111111"), -- 19 (fails: pc)
      -- ("2B67"            , "F4D0"            , '0', "0000"            , '0', "03E8"           , "000A"           , "FFFF"            )
         ("0010101101100111", "0000000000001110", '0', "----------------", '0', "000001111101000", "000000000001010", "1111111111111111"), -- 20 (fails: pc)
      -- ("2B67"            , "000E"            , '0', "0000"            , '0', "03E8"           , "000A"           , "FFFF"            )
         ("0010101101100111", "0000000000001110", '0', "----------------", '0', "000000000001110", "000000000001011", "1111111111111111"), -- 21 (fails: pc)
      -- ("2B67"            , "000E"            , '0', "0000"            , '0', "000E"           , "000B"           , "FFFF"            )
         ("0010101101100111", "1110001100000100", '0', "----------------", '0', "000000000001110", "000000000001011", "1111111111111111"), -- 22 (fails: pc)
      -- ("2B67"            , "E304"            , '0', "0000"            , '0', "000E"           , "000B"           , "FFFF"            )
         ("0010101101100111", "1110001100000100", '0', "----------------", '0', "000000000001110", "000000000001110", "1111111111111111"), -- 23 (fails: pc)
      -- ("2B67"            , "E304"            , '0', "0000"            , '0', "000E"           , "000E"           , "FFFF"            )
         ("0010101101100111", "0000001111100111", '0', "----------------", '0', "000000000001110", "000000000001110", "1111111111111111"), -- 24 (fails: pc)
      -- ("2B67"            , "03E7"            , '0', "0000"            , '0', "000E"           , "000E"           , "FFFF"            )
         ("0010101101100111", "0000001111100111", '0', "----------------", '0', "000001111100111", "000000000001111", "1111111111111111"), -- 25 (fails: pc)
      -- ("2B67"            , "03E7"            , '0', "0000"            , '0', "03E7"           , "000F"           , "FFFF"            )
         ("0010101101100111", "1110110111100000", '0', "----------------", '0', "000001111100111", "000000000001111", "1111111111111111"), -- 26 (fails: pc)
      -- ("2B67"            , "EDE0"            , '0', "0000"            , '0', "03E7"           , "000F"           , "FFFF"            )
         ("0010101101100111", "1110110111100000", '0', "----------------", '0', "000001111101000", "000000000010000", "1111111111111111"), -- 27 (fails: pc)
      -- ("2B67"            , "EDE0"            , '0', "0000"            , '0', "03E8"           , "0010"           , "FFFF"            )
         ("0010101101100111", "1110001100001000", '0', "1111111111111111", '1', "000001111101000", "000000000010000", "1111111111111111"), -- 28 (fails: addressM cpu tb)
      -- ("2B67"            , "E308"            , '0', "FFFF"            , '1', "03E8"           , "0010"           , "FFFF"            )
         ("0010101101100111", "1110001100001000", '0', "1111111111111111", '1', "000001111101000", "000000000010001", "1111111111111111"), -- 29 (fails: addressM cpu pc)
      -- ("2B67"            , "E308"            , '0', "FFFF"            , '1', "03E8"           , "0011"           , "FFFF"            )
         ("0010101101100111", "0000000000010101", '0', "----------------", '0', "000001111101000", "000000000010001", "1111111111111111"), -- 30 (fails: addressM pc)
      -- ("2B67"            , "0015"            , '0', "0000"            , '0', "03E8"           , "0011"           , "FFFF"            )
         ("0010101101100111", "0000000000010101", '0', "----------------", '0', "000000000010101", "000000000010010", "1111111111111111"), -- 31 (fails: pc)
      -- ("2B67"            , "0015"            , '0', "0000"            , '0', "0015"           , "0012"           , "FFFF"            )
         ("0010101101100111", "1110011111000010", '0', "----------------", '0', "000000000010101", "000000000010010", "1111111111111111"), -- 32 (fails: pc)
      -- ("2B67"            , "E7C2"            , '0', "0000"            , '0', "0015"           , "0012"           , "FFFF"            )
         ("0010101101100111", "1110011111000010", '0', "----------------", '0', "000000000010101", "000000000010101", "1111111111111111"), -- 33 (fails: pc)
      -- ("2B67"            , "E7C2"            , '0', "0000"            , '0', "0015"           , "0015"           , "FFFF"            )
         ("0010101101100111", "0000000000000010", '0', "----------------", '0', "000000000010101", "000000000010101", "1111111111111111"), -- 34 (fails: pc)
      -- ("2B67"            , "0002"            , '0', "0000"            , '0', "0015"           , "0015"           , "FFFF"            )
         ("0010101101100111", "0000000000000010", '0', "----------------", '0', "000000000000010", "000000000010110", "1111111111111111"), -- 35 (fails: pc)
      -- ("2B67"            , "0002"            , '0', "0000"            , '0', "0002"           , "0016"           , "FFFF"            )
         ("0010101101100111", "1110000010010000", '0', "----------------", '0', "000000000000010", "000000000010110", "0000000000000001"), -- 36 (fails: pc)
      -- ("2B67"            , "E090"            , '0', "0000"            , '0', "0002"           , "0016"           , "0001"            )
         ("0010101101100111", "1110000010010000", '0', "----------------", '0', "000000000000010", "000000000010111", "0000000000000001"), -- 37 (fails: pc)
      -- ("2B67"            , "E090"            , '0', "0000"            , '0', "0002"           , "0017"           , "0001"            )
         ("0010101101100111", "0000001111101000", '0', "----------------", '0', "000000000000010", "000000000010111", "0000000000000001"), -- 38 (fails: pc)
      -- ("2B67"            , "03E8"            , '0', "0000"            , '0', "0002"           , "0017"           , "0001"            )
         ("0010101101100111", "0000001111101000", '0', "----------------", '0', "000001111101000", "000000000011000", "0000000000000001"), -- 39 (fails: pc)
      -- ("2B67"            , "03E8"            , '0', "0000"            , '0', "03E8"           , "0018"           , "0001"            )
         ("0010101101100111", "1110111010010000", '0', "----------------", '0', "000001111101000", "000000000011000", "1111111111111111"), -- 40 (fails: pc)
      -- ("2B67"            , "EE90"            , '0', "0000"            , '0', "03E8"           , "0018"           , "FFFF"            )
         ("0010101101100111", "1110111010010000", '0', "----------------", '0', "000001111101000", "000000000011001", "1111111111111111"), -- 41 (fails: pc)
      -- ("2B67"            , "EE90"            , '0', "0000"            , '0', "03E8"           , "0019"           , "FFFF"            )
         ("0010101101100111", "1110001100000001", '0', "----------------", '0', "000001111101000", "000000000011001", "1111111111111111"), -- 42 (fails: pc)
      -- ("2B67"            , "E301"            , '0', "0000"            , '0', "03E8"           , "0019"           , "FFFF"            )
         ("0010101101100111", "1110001100000001", '0', "----------------", '0', "000001111101000", "000000000011010", "1111111111111111"), -- 43 (fails: pc)
      -- ("2B67"            , "E301"            , '0', "0000"            , '0', "03E8"           , "001A"           , "FFFF"            )
         ("0010101101100111", "1110001100000010", '0', "----------------", '0', "000001111101000", "000000000011010", "1111111111111111"), -- 44 (fails: pc)
      -- ("2B67"            , "E302"            , '0', "0000"            , '0', "03E8"           , "001A"           , "FFFF"            )
         ("0010101101100111", "1110001100000010", '0', "----------------", '0', "000001111101000", "000000000011011", "1111111111111111"), -- 45 (fails: pc)
      -- ("2B67"            , "E302"            , '0', "0000"            , '0', "03E8"           , "001B"           , "FFFF"            )
         ("0010101101100111", "1110001100000011", '0', "----------------", '0', "000001111101000", "000000000011011", "1111111111111111"), -- 46 (fails: pc)
      -- ("2B67"            , "E303"            , '0', "0000"            , '0', "03E8"           , "001B"           , "FFFF"            )
         ("0010101101100111", "1110001100000011", '0', "----------------", '0', "000001111101000", "000000000011100", "1111111111111111"), -- 47 (fails: pc)
      -- ("2B67"            , "E303"            , '0', "0000"            , '0', "03E8"           , "001C"           , "FFFF"            )
         ("0010101101100111", "1110001100000100", '0', "----------------", '0', "000001111101000", "000000000011100", "1111111111111111"), -- 48 (fails: pc)
      -- ("2B67"            , "E304"            , '0', "0000"            , '0', "03E8"           , "001C"           , "FFFF"            )
         ("0010101101100111", "1110001100000100", '0', "----------------", '0', "000001111101000", "000001111101000", "1111111111111111"), -- 49 (fails: pc)
      -- ("2B67"            , "E304"            , '0', "0000"            , '0', "03E8"           , "03E8"           , "FFFF"            )
         ("0010101101100111", "1110001100000101", '0', "----------------", '0', "000001111101000", "000001111101000", "1111111111111111"), -- 50 (fails: pc)
      -- ("2B67"            , "E305"            , '0', "0000"            , '0', "03E8"           , "03E8"           , "FFFF"            )
         ("0010101101100111", "1110001100000101", '0', "----------------", '0', "000001111101000", "000001111101000", "1111111111111111"), -- 51 (fails: pc)
      -- ("2B67"            , "E305"            , '0', "0000"            , '0', "03E8"           , "03E8"           , "FFFF"            )
         ("0010101101100111", "1110001100000110", '0', "----------------", '0', "000001111101000", "000001111101000", "1111111111111111"), -- 52 (fails: pc)
      -- ("2B67"            , "E306"            , '0', "0000"            , '0', "03E8"           , "03E8"           , "FFFF"            )
         ("0010101101100111", "1110001100000110", '0', "----------------", '0', "000001111101000", "000001111101000", "1111111111111111"), -- 53 (fails: pc)
      -- ("2B67"            , "E306"            , '0', "0000"            , '0', "03E8"           , "03E8"           , "FFFF"            )
         ("0010101101100111", "1110001100000111", '0', "----------------", '0', "000001111101000", "000001111101000", "1111111111111111"), -- 54 (fails: pc)
      -- ("2B67"            , "E307"            , '0', "0000"            , '0', "03E8"           , "03E8"           , "FFFF"            )
         ("0010101101100111", "1110001100000111", '0', "----------------", '0', "000001111101000", "000001111101000", "1111111111111111"), -- 55 (fails: pc)
      -- ("2B67"            , "E307"            , '0', "0000"            , '0', "03E8"           , "03E8"           , "FFFF"            )
         ("0010101101100111", "1110101010010000", '0', "----------------", '0', "000001111101000", "000001111101000", "0000000000000000"), -- 56 (fails: pc)
      -- ("2B67"            , "EA90"            , '0', "0000"            , '0', "03E8"           , "03E8"           , "0000"            )
         ("0010101101100111", "1110101010010000", '0', "----------------", '0', "000001111101000", "000001111101001", "0000000000000000"), -- 57 (fails: pc)
      -- ("2B67"            , "EA90"            , '0', "0000"            , '0', "03E8"           , "03E9"           , "0000"            )
         ("0010101101100111", "1110001100000001", '0', "----------------", '0', "000001111101000", "000001111101001", "0000000000000000"), -- 58 (fails: pc)
      -- ("2B67"            , "E301"            , '0', "0000"            , '0', "03E8"           , "03E9"           , "0000"            )
         ("0010101101100111", "1110001100000001", '0', "----------------", '0', "000001111101000", "000001111101010", "0000000000000000"), -- 59 (fails: pc)
      -- ("2B67"            , "E301"            , '0', "0000"            , '0', "03E8"           , "03EA"           , "0000"            )
         ("0010101101100111", "1110001100000010", '0', "----------------", '0', "000001111101000", "000001111101010", "0000000000000000"), -- 60 (fails: pc)
      -- ("2B67"            , "E302"            , '0', "0000"            , '0', "03E8"           , "03EA"           , "0000"            )
         ("0010101101100111", "1110001100000010", '0', "----------------", '0', "000001111101000", "000001111101000", "0000000000000000"), -- 61 (fails: pc)
      -- ("2B67"            , "E302"            , '0', "0000"            , '0', "03E8"           , "03E8"           , "0000"            )
         ("0010101101100111", "1110001100000011", '0', "----------------", '0', "000001111101000", "000001111101000", "0000000000000000"), -- 62 (fails: pc)
      -- ("2B67"            , "E303"            , '0', "0000"            , '0', "03E8"           , "03E8"           , "0000"            )
         ("0010101101100111", "1110001100000011", '0', "----------------", '0', "000001111101000", "000001111101000", "0000000000000000"), -- 63 (fails: pc)
      -- ("2B67"            , "E303"            , '0', "0000"            , '0', "03E8"           , "03E8"           , "0000"            )
         ("0010101101100111", "1110001100000100", '0', "----------------", '0', "000001111101000", "000001111101000", "0000000000000000"), -- 64 (fails: pc)
      -- ("2B67"            , "E304"            , '0', "0000"            , '0', "03E8"           , "03E8"           , "0000"            )
         ("0010101101100111", "1110001100000100", '0', "----------------", '0', "000001111101000", "000001111101001", "0000000000000000"), -- 65 (fails: pc)
      -- ("2B67"            , "E304"            , '0', "0000"            , '0', "03E8"           , "03E9"           , "0000"            )
         ("0010101101100111", "1110001100000101", '0', "----------------", '0', "000001111101000", "000001111101001", "0000000000000000"), -- 66 (fails: pc)
      -- ("2B67"            , "E305"            , '0', "0000"            , '0', "03E8"           , "03E9"           , "0000"            )
         ("0010101101100111", "1110001100000101", '0', "----------------", '0', "000001111101000", "000001111101010", "0000000000000000"), -- 67 (fails: pc)
      -- ("2B67"            , "E305"            , '0', "0000"            , '0', "03E8"           , "03EA"           , "0000"            )
         ("0010101101100111", "1110001100000110", '0', "----------------", '0', "000001111101000", "000001111101010", "0000000000000000"), -- 68 (fails: pc)
      -- ("2B67"            , "E306"            , '0', "0000"            , '0', "03E8"           , "03EA"           , "0000"            )
         ("0010101101100111", "1110001100000110", '0', "----------------", '0', "000001111101000", "000001111101000", "0000000000000000"), -- 69 (fails: pc)
      -- ("2B67"            , "E306"            , '0', "0000"            , '0', "03E8"           , "03E8"           , "0000"            )
         ("0010101101100111", "1110001100000111", '0', "----------------", '0', "000001111101000", "000001111101000", "0000000000000000"), -- 70 (fails: pc)
      -- ("2B67"            , "E307"            , '0', "0000"            , '0', "03E8"           , "03E8"           , "0000"            )
         ("0010101101100111", "1110001100000111", '0', "----------------", '0', "000001111101000", "000001111101000", "0000000000000000"), -- 71 (fails: pc)
      -- ("2B67"            , "E307"            , '0', "0000"            , '0', "03E8"           , "03E8"           , "0000"            )
         ("0010101101100111", "1110111111010000", '0', "----------------", '0', "000001111101000", "000001111101000", "0000000000000001"), -- 72 (fails: pc)
      -- ("2B67"            , "EFD0"            , '0', "0000"            , '0', "03E8"           , "03E8"           , "0001"            )
         ("0010101101100111", "1110111111010000", '0', "----------------", '0', "000001111101000", "000001111101001", "0000000000000001"), -- 73 (fails: pc)
      -- ("2B67"            , "EFD0"            , '0', "0000"            , '0', "03E8"           , "03E9"           , "0001"            )
         ("0010101101100111", "1110001100000001", '0', "----------------", '0', "000001111101000", "000001111101001", "0000000000000001"), -- 74 (fails: pc)
      -- ("2B67"            , "E301"            , '0', "0000"            , '0', "03E8"           , "03E9"           , "0001"            )
         ("0010101101100111", "1110001100000001", '0', "----------------", '0', "000001111101000", "000001111101000", "0000000000000001"), -- 75 (fails: pc)
      -- ("2B67"            , "E301"            , '0', "0000"            , '0', "03E8"           , "03E8"           , "0001"            )
         ("0010101101100111", "1110001100000010", '0', "----------------", '0', "000001111101000", "000001111101000", "0000000000000001"), -- 76 (fails: pc)
      -- ("2B67"            , "E302"            , '0', "0000"            , '0', "03E8"           , "03E8"           , "0001"            )
         ("0010101101100111", "1110001100000010", '0', "----------------", '0', "000001111101000", "000001111101001", "0000000000000001"), -- 77 (fails: pc)
      -- ("2B67"            , "E302"            , '0', "0000"            , '0', "03E8"           , "03E9"           , "0001"            )
         ("0010101101100111", "1110001100000011", '0', "----------------", '0', "000001111101000", "000001111101001", "0000000000000001"), -- 78 (fails: pc)
      -- ("2B67"            , "E303"            , '0', "0000"            , '0', "03E8"           , "03E9"           , "0001"            )
         ("0010101101100111", "1110001100000011", '0', "----------------", '0', "000001111101000", "000001111101000", "0000000000000001"), -- 79 (fails: pc)
      -- ("2B67"            , "E303"            , '0', "0000"            , '0', "03E8"           , "03E8"           , "0001"            )
         ("0010101101100111", "1110001100000100", '0', "----------------", '0', "000001111101000", "000001111101000", "0000000000000001"), -- 80 (fails: pc)
      -- ("2B67"            , "E304"            , '0', "0000"            , '0', "03E8"           , "03E8"           , "0001"            )
         ("0010101101100111", "1110001100000100", '0', "----------------", '0', "000001111101000", "000001111101001", "0000000000000001"), -- 81 (fails: pc)
      -- ("2B67"            , "E304"            , '0', "0000"            , '0', "03E8"           , "03E9"           , "0001"            )
         ("0010101101100111", "1110001100000101", '0', "----------------", '0', "000001111101000", "000001111101001", "0000000000000001"), -- 82 (fails: pc)
      -- ("2B67"            , "E305"            , '0', "0000"            , '0', "03E8"           , "03E9"           , "0001"            )
         ("0010101101100111", "1110001100000101", '0', "----------------", '0', "000001111101000", "000001111101000", "0000000000000001"), -- 83 (fails: pc)
      -- ("2B67"            , "E305"            , '0', "0000"            , '0', "03E8"           , "03E8"           , "0001"            )
         ("0010101101100111", "1110001100000110", '0', "----------------", '0', "000001111101000", "000001111101000", "0000000000000001"), -- 84 (fails: pc)
      -- ("2B67"            , "E306"            , '0', "0000"            , '0', "03E8"           , "03E8"           , "0001"            )
         ("0010101101100111", "1110001100000110", '0', "----------------", '0', "000001111101000", "000001111101001", "0000000000000001"), -- 85 (fails: pc)
      -- ("2B67"            , "E306"            , '0', "0000"            , '0', "03E8"           , "03E9"           , "0001"            )
         ("0010101101100111", "1110001100000111", '0', "----------------", '0', "000001111101000", "000001111101001", "0000000000000001"), -- 86 (fails: pc)
      -- ("2B67"            , "E307"            , '0', "0000"            , '0', "03E8"           , "03E9"           , "0001"            )
         ("0010101101100111", "1110001100000111", '0', "----------------", '0', "000001111101000", "000001111101000", "0000000000000001"), -- 87 (fails: pc)
      -- ("2B67"            , "E307"            , '0', "0000"            , '0', "03E8"           , "03E8"           , "0001"            )
         ("0010101101100111", "1110001100000111", '1', "----------------", '0', "000001111101000", "000001111101000", "0000000000000001"), -- 88 (fails: pc)
      -- ("2B67"            , "E307"            , '1', "0000"            , '0', "03E8"           , "03E8"           , "0001"            )
         ("0010101101100111", "1110001100000111", '1', "----------------", '0', "000001111101000", "000000000000000", "0000000000000001"), -- 89 (fails: pc)
      -- ("2B67"            , "E307"            , '1', "0000"            , '0', "03E8"           , "0000"           , "0001"            )
         ("0010101101100111", "0111111111111111", '0', "----------------", '0', "000001111101000", "000000000000000", "0000000000000001"), -- 90 (fails: pc)
      -- ("2B67"            , "7FFF"            , '0', "0000"            , '0', "03E8"           , "0000"           , "0001"            )
         ("0010101101100111", "0111111111111111", '0', "----------------", '0', "111111111111111", "000000000000001", "0000000000000001")); -- 91 (fails: pc)
      -- ("2B67"            , "7FFF"            , '0', "0000"            , '0', "7FFF"           , "0001"           , "0001"            )
         
   begin
      --  Check each pattern.
      for i in patterns'range loop
         --  Set the inputs.
         inM <= patterns(i).inM;
         instruction <= patterns(i).instruction;
         reset <= patterns(i).reset;

         -- Wait for the results
         wait for 0.25 ns;

         --  Check the outputs.
         if (patterns(i).outM /= "----------------") then
           assert outM = patterns(i).outM
             report "bad cpu output" severity error;
         end if;
         assert writeM = patterns(i).writeM
           report "bad writeM output bit" severity error;
         assert addressM = patterns(i).addressM
           report "bad addressM output" severity error;
         assert pcOut = patterns(i).pcOut
           report "bad pc output" severity error;

         -- Wait the rest of the cycle
         wait for 0.75 ns;
      end loop;

      -- End the clock
      finish <= '1';

      assert false report "end of test" severity note;
      --  Wait forever; this will finish the simulation.
      wait;
   end process;
end cpu_tb_arch;
