library IEEE;
use IEEE.std_logic_1164.all;

--  A testbench has no ports.
entity ram64_tb is
end ram64_tb;

architecture ram64_tb_arch of ram64_tb is
   --  Declaration of the component that will be instantiated.
   component ram64
     port (d       : in std_logic_vector(15 downto 0);
           load    : in std_logic;
           address : in std_logic_vector(5 downto 0);
           clk     : in std_logic;
           cout    : out std_logic_vector(15 downto 0));
   end component;
   -- Declaration of the clock
   component Clock
     port (finish : in std_logic;
           cout   : out std_logic);
   end component;
   
   --  Specifies which entity is bound with the component.
   for ram64_0: ram64 use entity work.ram64;
   signal d, cout : std_logic_vector(15 downto 0);
   signal address : std_logic_vector(5 downto 0);
   signal load, finish, clk : std_logic;
begin
  --  Component instantiation.
  OSC_CLK: Clock port map (finish, clk);
  ram64_0: ram64 port map (d, load, address, clk, cout);

   --  This process does the real job.
   process
      type pattern_type is record
         --  The inputs of the ram64.
        d       : std_logic_vector(15 downto 0);
        load    : std_logic;
        address : std_logic_vector(5 downto 0);
        --  The output of the ram64.
        cout    : std_logic_vector(15 downto 0);
      end record;
      --  The patterns to apply.
      type pattern_array is array (natural range <>) of pattern_type;
      constant patterns : pattern_array :=
        (("0000000000000000", '0', "000000", "0000000000000000"),
         ("0000000000000000", '0', "000000", "0000000000000000"),
         ("0000000000000000", '1', "000000", "0000000000000000"),
         ("0000000000000000", '1', "000000", "0000000000000000"),
         ("0000010100100001", '0', "000000", "0000000000000000"),
         ("0000010100100001", '0', "000000", "0000000000000000"),
         ("0000010100100001", '1', "001101", "0000000000000000"),
         ("0000010100100001", '1', "001101", "0000010100100001"),
         ("0000010100100001", '0', "000000", "0000000000000000"),
         ("0000010100100001", '0', "000000", "0000000000000000"),
         ("0001001010001011", '0', "101111", "0000000000000000"),
         ("0001001010001011", '0', "101111", "0000000000000000"),
         ("0001001010001011", '1', "101111", "0000000000000000"),
         ("0001001010001011", '1', "101111", "0001001010001011"),
         ("0001001010001011", '0', "101111", "0001001010001011"),
         ("0001001010001011", '0', "101111", "0001001010001011"),
         ("0001001010001011", '0', "001101", "0000010100100001"),
         ("0001100011011011", '0', "001101", "0000010100100001"),
         ("0001100011011011", '0', "001101", "0000010100100001"),
         ("0001100011011011", '1', "111111", "0000000000000000"),
         ("0001100011011011", '1', "111111", "0001100011011011"),
         ("0001100011011011", '0', "111111", "0001100011011011"),
         ("0001100011011011", '0', "111111", "0001100011011011"),
         ("0001100011011011", '0', "101111", "0001001010001011"),
         ("0001100011011011", '0', "111111", "0001100011011011"),
         ("0001100011011011", '0', "101000", "0000000000000000"),
         ("0001100011011011", '0', "101000", "0000000000000000"),
         ("0001100011011011", '0', "101001", "0000000000000000"),
         ("0001100011011011", '0', "101010", "0000000000000000"),
         ("0001100011011011", '0', "101011", "0000000000000000"),
         ("0001100011011011", '0', "101100", "0000000000000000"),
         ("0001100011011011", '0', "101101", "0000000000000000"),
         ("0001100011011011", '0', "101110", "0000000000000000"),
         ("0001100011011011", '0', "101111", "0001001010001011"),
         ("0101010101010101", '1', "101000", "0000000000000000"),
         ("0101010101010101", '1', "101000", "0101010101010101"),
         ("0101010101010101", '1', "101001", "0000000000000000"),
         ("0101010101010101", '1', "101001", "0101010101010101"),
         ("0101010101010101", '1', "101010", "0000000000000000"),
         ("0101010101010101", '1', "101010", "0101010101010101"),
         ("0101010101010101", '1', "101011", "0000000000000000"),
         ("0101010101010101", '1', "101011", "0101010101010101"),
         ("0101010101010101", '1', "101100", "0000000000000000"),
         ("0101010101010101", '1', "101100", "0101010101010101"),
         ("0101010101010101", '1', "101101", "0000000000000000"),
         ("0101010101010101", '1', "101101", "0101010101010101"),
         ("0101010101010101", '1', "101110", "0000000000000000"),
         ("0101010101010101", '1', "101110", "0101010101010101"),
         ("0101010101010101", '1', "101111", "0001001010001011"),
         ("0101010101010101", '1', "101111", "0101010101010101"),
         ("0101010101010101", '0', "101000", "0101010101010101"),
         ("0101010101010101", '0', "101000", "0101010101010101"),
         ("0101010101010101", '0', "101001", "0101010101010101"),
         ("0101010101010101", '0', "101010", "0101010101010101"),
         ("0101010101010101", '0', "101011", "0101010101010101"),
         ("0101010101010101", '0', "101100", "0101010101010101"),
         ("0101010101010101", '0', "101101", "0101010101010101"),
         ("0101010101010101", '0', "101110", "0101010101010101"),
         ("0101010101010101", '0', "101111", "0101010101010101"),
         ("0101010101010110", '1', "101000", "0101010101010101"),
         ("0101010101010110", '1', "101000", "0101010101010110"),
         ("0101010101010110", '0', "101000", "0101010101010110"),
         ("0101010101010110", '0', "101000", "0101010101010110"),
         ("0101010101010110", '0', "101001", "0101010101010101"),
         ("0101010101010110", '0', "101010", "0101010101010101"),
         ("0101010101010110", '0', "101011", "0101010101010101"),
         ("0101010101010110", '0', "101100", "0101010101010101"),
         ("0101010101010110", '0', "101101", "0101010101010101"),
         ("0101010101010110", '0', "101110", "0101010101010101"),
         ("0101010101010110", '0', "101111", "0101010101010101"),
         ("0101010101010101", '1', "101000", "0101010101010110"),
         ("0101010101010101", '1', "101000", "0101010101010101"),
         ("0101010101010110", '1', "101001", "0101010101010101"),
         ("0101010101010110", '1', "101001", "0101010101010110"),
         ("0101010101010110", '0', "101000", "0101010101010101"),
         ("0101010101010110", '0', "101000", "0101010101010101"),
         ("0101010101010110", '0', "101001", "0101010101010110"),
         ("0101010101010110", '0', "101010", "0101010101010101"),
         ("0101010101010110", '0', "101011", "0101010101010101"),
         ("0101010101010110", '0', "101100", "0101010101010101"),
         ("0101010101010110", '0', "101101", "0101010101010101"),
         ("0101010101010110", '0', "101110", "0101010101010101"),
         ("0101010101010110", '0', "101111", "0101010101010101"),
         ("0101010101010101", '1', "101001", "0101010101010110"),
         ("0101010101010101", '1', "101001", "0101010101010101"),
         ("0101010101010110", '1', "101010", "0101010101010101"),
         ("0101010101010110", '1', "101010", "0101010101010110"),
         ("0101010101010110", '0', "101000", "0101010101010101"),
         ("0101010101010110", '0', "101000", "0101010101010101"),
         ("0101010101010110", '0', "101001", "0101010101010101"),
         ("0101010101010110", '0', "101010", "0101010101010110"),
         ("0101010101010110", '0', "101011", "0101010101010101"),
         ("0101010101010110", '0', "101100", "0101010101010101"),
         ("0101010101010110", '0', "101101", "0101010101010101"),
         ("0101010101010110", '0', "101110", "0101010101010101"),
         ("0101010101010110", '0', "101111", "0101010101010101"),
         ("0101010101010101", '1', "101010", "0101010101010110"),
         ("0101010101010101", '1', "101010", "0101010101010101"),
         ("0101010101010110", '1', "101011", "0101010101010101"),
         ("0101010101010110", '1', "101011", "0101010101010110"),
         ("0101010101010110", '0', "101000", "0101010101010101"),
         ("0101010101010110", '0', "101000", "0101010101010101"),
         ("0101010101010110", '0', "101001", "0101010101010101"),
         ("0101010101010110", '0', "101010", "0101010101010101"),
         ("0101010101010110", '0', "101011", "0101010101010110"),
         ("0101010101010110", '0', "101100", "0101010101010101"),
         ("0101010101010110", '0', "101101", "0101010101010101"),
         ("0101010101010110", '0', "101110", "0101010101010101"),
         ("0101010101010110", '0', "101111", "0101010101010101"),
         ("0101010101010101", '1', "101011", "0101010101010110"),
         ("0101010101010101", '1', "101011", "0101010101010101"),
         ("0101010101010110", '1', "101100", "0101010101010101"),
         ("0101010101010110", '1', "101100", "0101010101010110"),
         ("0101010101010110", '0', "101000", "0101010101010101"),
         ("0101010101010110", '0', "101000", "0101010101010101"),
         ("0101010101010110", '0', "101001", "0101010101010101"),
         ("0101010101010110", '0', "101010", "0101010101010101"),
         ("0101010101010110", '0', "101011", "0101010101010101"),
         ("0101010101010110", '0', "101100", "0101010101010110"),
         ("0101010101010110", '0', "101101", "0101010101010101"),
         ("0101010101010110", '0', "101110", "0101010101010101"),
         ("0101010101010110", '0', "101111", "0101010101010101"),
         ("0101010101010101", '1', "101100", "0101010101010110"),
         ("0101010101010101", '1', "101100", "0101010101010101"),
         ("0101010101010110", '1', "101101", "0101010101010101"),
         ("0101010101010110", '1', "101101", "0101010101010110"),
         ("0101010101010110", '0', "101000", "0101010101010101"),
         ("0101010101010110", '0', "101000", "0101010101010101"),
         ("0101010101010110", '0', "101001", "0101010101010101"),
         ("0101010101010110", '0', "101010", "0101010101010101"),
         ("0101010101010110", '0', "101011", "0101010101010101"),
         ("0101010101010110", '0', "101100", "0101010101010101"),
         ("0101010101010110", '0', "101101", "0101010101010110"),
         ("0101010101010110", '0', "101110", "0101010101010101"),
         ("0101010101010110", '0', "101111", "0101010101010101"),
         ("0101010101010101", '1', "101101", "0101010101010110"),
         ("0101010101010101", '1', "101101", "0101010101010101"),
         ("0101010101010110", '1', "101110", "0101010101010101"),
         ("0101010101010110", '1', "101110", "0101010101010110"),
         ("0101010101010110", '0', "101000", "0101010101010101"),
         ("0101010101010110", '0', "101000", "0101010101010101"),
         ("0101010101010110", '0', "101001", "0101010101010101"),
         ("0101010101010110", '0', "101010", "0101010101010101"),
         ("0101010101010110", '0', "101011", "0101010101010101"),
         ("0101010101010110", '0', "101100", "0101010101010101"),
         ("0101010101010110", '0', "101101", "0101010101010101"),
         ("0101010101010110", '0', "101110", "0101010101010110"),
         ("0101010101010110", '0', "101111", "0101010101010101"),
         ("0101010101010101", '1', "101110", "0101010101010110"),
         ("0101010101010101", '1', "101110", "0101010101010101"),
         ("0101010101010110", '1', "101111", "0101010101010101"),
         ("0101010101010110", '1', "101111", "0101010101010110"),
         ("0101010101010110", '0', "101000", "0101010101010101"),
         ("0101010101010110", '0', "101000", "0101010101010101"),
         ("0101010101010110", '0', "101001", "0101010101010101"),
         ("0101010101010110", '0', "101010", "0101010101010101"),
         ("0101010101010110", '0', "101011", "0101010101010101"),
         ("0101010101010110", '0', "101100", "0101010101010101"),
         ("0101010101010110", '0', "101101", "0101010101010101"),
         ("0101010101010110", '0', "101110", "0101010101010101"),
         ("0101010101010110", '0', "101111", "0101010101010110"),
         ("0101010101010101", '1', "101111", "0101010101010110"),
         ("0101010101010101", '1', "101111", "0101010101010101"),
         ("0101010101010101", '0', "101000", "0101010101010101"),
         ("0101010101010101", '0', "101000", "0101010101010101"),
         ("0101010101010101", '0', "101001", "0101010101010101"),
         ("0101010101010101", '0', "101010", "0101010101010101"),
         ("0101010101010101", '0', "101011", "0101010101010101"),
         ("0101010101010101", '0', "101100", "0101010101010101"),
         ("0101010101010101", '0', "101101", "0101010101010101"),
         ("0101010101010101", '0', "101110", "0101010101010101"),
         ("0101010101010101", '0', "101111", "0101010101010101"),
         ("0101010101010101", '0', "000101", "0000000000000000"),
         ("0101010101010101", '0', "000101", "0000000000000000"),
         ("0101010101010101", '0', "001101", "0000010100100001"),
         ("0101010101010101", '0', "010101", "0000000000000000"),
         ("0101010101010101", '0', "011101", "0000000000000000"),
         ("0101010101010101", '0', "100101", "0000000000000000"),
         ("0101010101010101", '0', "101101", "0101010101010101"),
         ("0101010101010101", '0', "110101", "0000000000000000"),
         ("0101010101010101", '0', "111101", "0000000000000000"),
         ("0101010101010101", '1', "000101", "0000000000000000"),
         ("0101010101010101", '1', "000101", "0101010101010101"),
         ("0101010101010101", '1', "001101", "0000010100100001"),
         ("0101010101010101", '1', "001101", "0101010101010101"),
         ("0101010101010101", '1', "010101", "0000000000000000"),
         ("0101010101010101", '1', "010101", "0101010101010101"),
         ("0101010101010101", '1', "011101", "0000000000000000"),
         ("0101010101010101", '1', "011101", "0101010101010101"),
         ("0101010101010101", '1', "100101", "0000000000000000"),
         ("0101010101010101", '1', "100101", "0101010101010101"),
         ("0101010101010101", '1', "101101", "0101010101010101"),
         ("0101010101010101", '1', "101101", "0101010101010101"),
         ("0101010101010101", '1', "110101", "0000000000000000"),
         ("0101010101010101", '1', "110101", "0101010101010101"),
         ("0101010101010101", '1', "111101", "0000000000000000"),
         ("0101010101010101", '1', "111101", "0101010101010101"),
         ("0101010101010101", '0', "000101", "0101010101010101"),
         ("0101010101010101", '0', "000101", "0101010101010101"),
         ("0101010101010101", '0', "001101", "0101010101010101"),
         ("0101010101010101", '0', "010101", "0101010101010101"),
         ("0101010101010101", '0', "011101", "0101010101010101"),
         ("0101010101010101", '0', "100101", "0101010101010101"),
         ("0101010101010101", '0', "101101", "0101010101010101"),
         ("0101010101010101", '0', "110101", "0101010101010101"),
         ("0101010101010101", '0', "111101", "0101010101010101"),
         ("0101010101010110", '1', "000101", "0101010101010101"),
         ("0101010101010110", '1', "000101", "0101010101010110"),
         ("0101010101010110", '0', "000101", "0101010101010110"),
         ("0101010101010110", '0', "000101", "0101010101010110"),
         ("0101010101010110", '0', "001101", "0101010101010101"),
         ("0101010101010110", '0', "010101", "0101010101010101"),
         ("0101010101010110", '0', "011101", "0101010101010101"),
         ("0101010101010110", '0', "100101", "0101010101010101"),
         ("0101010101010110", '0', "101101", "0101010101010101"),
         ("0101010101010110", '0', "110101", "0101010101010101"),
         ("0101010101010110", '0', "111101", "0101010101010101"),
         ("0101010101010101", '1', "000101", "0101010101010110"),
         ("0101010101010101", '1', "000101", "0101010101010101"),
         ("0101010101010110", '1', "001101", "0101010101010101"),
         ("0101010101010110", '1', "001101", "0101010101010110"),
         ("0101010101010110", '0', "000101", "0101010101010101"),
         ("0101010101010110", '0', "000101", "0101010101010101"),
         ("0101010101010110", '0', "001101", "0101010101010110"),
         ("0101010101010110", '0', "010101", "0101010101010101"),
         ("0101010101010110", '0', "011101", "0101010101010101"),
         ("0101010101010110", '0', "100101", "0101010101010101"),
         ("0101010101010110", '0', "101101", "0101010101010101"),
         ("0101010101010110", '0', "110101", "0101010101010101"),
         ("0101010101010110", '0', "111101", "0101010101010101"),
         ("0101010101010101", '1', "001101", "0101010101010110"),
         ("0101010101010101", '1', "001101", "0101010101010101"),
         ("0101010101010110", '1', "010101", "0101010101010101"),
         ("0101010101010110", '1', "010101", "0101010101010110"),
         ("0101010101010110", '0', "000101", "0101010101010101"),
         ("0101010101010110", '0', "000101", "0101010101010101"),
         ("0101010101010110", '0', "001101", "0101010101010101"),
         ("0101010101010110", '0', "010101", "0101010101010110"),
         ("0101010101010110", '0', "011101", "0101010101010101"),
         ("0101010101010110", '0', "100101", "0101010101010101"),
         ("0101010101010110", '0', "101101", "0101010101010101"),
         ("0101010101010110", '0', "110101", "0101010101010101"),
         ("0101010101010110", '0', "111101", "0101010101010101"),
         ("0101010101010101", '1', "010101", "0101010101010110"),
         ("0101010101010101", '1', "010101", "0101010101010101"),
         ("0101010101010110", '1', "011101", "0101010101010101"),
         ("0101010101010110", '1', "011101", "0101010101010110"),
         ("0101010101010110", '0', "000101", "0101010101010101"),
         ("0101010101010110", '0', "000101", "0101010101010101"),
         ("0101010101010110", '0', "001101", "0101010101010101"),
         ("0101010101010110", '0', "010101", "0101010101010101"),
         ("0101010101010110", '0', "011101", "0101010101010110"),
         ("0101010101010110", '0', "100101", "0101010101010101"),
         ("0101010101010110", '0', "101101", "0101010101010101"),
         ("0101010101010110", '0', "110101", "0101010101010101"),
         ("0101010101010110", '0', "111101", "0101010101010101"),
         ("0101010101010101", '1', "011101", "0101010101010110"),
         ("0101010101010101", '1', "011101", "0101010101010101"),
         ("0101010101010110", '1', "100101", "0101010101010101"),
         ("0101010101010110", '1', "100101", "0101010101010110"),
         ("0101010101010110", '0', "000101", "0101010101010101"),
         ("0101010101010110", '0', "000101", "0101010101010101"),
         ("0101010101010110", '0', "001101", "0101010101010101"),
         ("0101010101010110", '0', "010101", "0101010101010101"),
         ("0101010101010110", '0', "011101", "0101010101010101"),
         ("0101010101010110", '0', "100101", "0101010101010110"),
         ("0101010101010110", '0', "101101", "0101010101010101"),
         ("0101010101010110", '0', "110101", "0101010101010101"),
         ("0101010101010110", '0', "111101", "0101010101010101"),
         ("0101010101010101", '1', "100101", "0101010101010110"),
         ("0101010101010101", '1', "100101", "0101010101010101"),
         ("0101010101010110", '1', "101101", "0101010101010101"),
         ("0101010101010110", '1', "101101", "0101010101010110"),
         ("0101010101010110", '0', "000101", "0101010101010101"),
         ("0101010101010110", '0', "000101", "0101010101010101"),
         ("0101010101010110", '0', "001101", "0101010101010101"),
         ("0101010101010110", '0', "010101", "0101010101010101"),
         ("0101010101010110", '0', "011101", "0101010101010101"),
         ("0101010101010110", '0', "100101", "0101010101010101"),
         ("0101010101010110", '0', "101101", "0101010101010110"),
         ("0101010101010110", '0', "110101", "0101010101010101"),
         ("0101010101010110", '0', "111101", "0101010101010101"),
         ("0101010101010101", '1', "101101", "0101010101010110"),
         ("0101010101010101", '1', "101101", "0101010101010101"),
         ("0101010101010110", '1', "110101", "0101010101010101"),
         ("0101010101010110", '1', "110101", "0101010101010110"),
         ("0101010101010110", '0', "000101", "0101010101010101"),
         ("0101010101010110", '0', "000101", "0101010101010101"),
         ("0101010101010110", '0', "001101", "0101010101010101"),
         ("0101010101010110", '0', "010101", "0101010101010101"),
         ("0101010101010110", '0', "011101", "0101010101010101"),
         ("0101010101010110", '0', "100101", "0101010101010101"),
         ("0101010101010110", '0', "101101", "0101010101010101"),
         ("0101010101010110", '0', "110101", "0101010101010110"),
         ("0101010101010110", '0', "111101", "0101010101010101"),
         ("0101010101010101", '1', "110101", "0101010101010110"),
         ("0101010101010101", '1', "110101", "0101010101010101"),
         ("0101010101010110", '1', "111101", "0101010101010101"),
         ("0101010101010110", '1', "111101", "0101010101010110"),
         ("0101010101010110", '0', "000101", "0101010101010101"),
         ("0101010101010110", '0', "000101", "0101010101010101"),
         ("0101010101010110", '0', "001101", "0101010101010101"),
         ("0101010101010110", '0', "010101", "0101010101010101"),
         ("0101010101010110", '0', "011101", "0101010101010101"),
         ("0101010101010110", '0', "100101", "0101010101010101"),
         ("0101010101010110", '0', "101101", "0101010101010101"),
         ("0101010101010110", '0', "110101", "0101010101010101"),
         ("0101010101010110", '0', "111101", "0101010101010110"),
         ("0101010101010101", '1', "111101", "0101010101010110"),
         ("0101010101010101", '1', "111101", "0101010101010101"),
         ("0101010101010101", '0', "000101", "0101010101010101"),
         ("0101010101010101", '0', "000101", "0101010101010101"),
         ("0101010101010101", '0', "001101", "0101010101010101"),
         ("0101010101010101", '0', "010101", "0101010101010101"),
         ("0101010101010101", '0', "011101", "0101010101010101"),
         ("0101010101010101", '0', "100101", "0101010101010101"),
         ("0101010101010101", '0', "101101", "0101010101010101"),
         ("0101010101010101", '0', "110101", "0101010101010101"),
         ("0101010101010101", '0', "111101", "0101010101010101"));
         
   begin
      --  Check each pattern.
      for i in patterns'range loop
         --  Set the inputs.
        d <= patterns(i).d;
        load <= patterns(i).load;
        address <= patterns(i).address;
        wait for 0.25 ns;
        --  Check the outputs.
        assert cout = patterns(i).cout
          report "bad data, memory problem" severity error;
        wait for 0.75 ns;
     end loop;
     -- End the clock
     finish <= '1';
     assert false report "end of test" severity note;
     --  Wait forever; this will finish the simulation.
     wait;
  end process;
end ram64_tb_arch;
